�� 
 m o d u l e   m e m   # (                                       / /    
         p a r a m e t e r     A D D R _ L E N     =   1 1       / /    
 )   (  
         i n p u t     c l k ,   r s t ,  
         i n p u t     [ A D D R _ L E N - 1 : 0 ]   a d d r ,   / /   m e m o r y   a d d r e s s  
         o u t p u t   r e g   [ 3 1 : 0 ]   r d _ d a t a ,     / /   d a t a   r e a d   o u t  
         i n p u t     w r _ r e q ,  
         i n p u t     [ 3 1 : 0 ]   w r _ d a t a               / /   d a t a   w r i t e   i n  
 ) ;  
 l o c a l p a r a m   M E M _ S I Z E   =   1 < < A D D R _ L E N ;  
 r e g   [ 3 1 : 0 ]   r a m _ c e l l   [ M E M _ S I Z E ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )  
                 r d _ d a t a   < =   0 ;  
         e l s e  
                 r d _ d a t a   < =   r a m _ c e l l [ a d d r ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k )  
         i f ( w r _ r e q )    
                 r a m _ c e l l [ a d d r ]   < =   w r _ d a t a ;  
  
 i n i t i a l   b e g i n  
         / /   d s t   m a t r i x   C  
         r a m _ c e l l [               0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 2 5 d 2 f 9 e ;  
         r a m _ c e l l [               1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 1 c b 0 d 8 4 ;  
         r a m _ c e l l [               2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 1 8 2 8 6 d e ;  
         r a m _ c e l l [               3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 0 d 2 7 c c c ;  
         r a m _ c e l l [               4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 9 c b a 0 b f ;  
         r a m _ c e l l [               5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 4 1 3 6 0 2 a ;  
         r a m _ c e l l [               6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 8 3 7 3 1 6 d ;  
         r a m _ c e l l [               7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 5 d 4 c f f d ;  
         r a m _ c e l l [               8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 5 6 7 a 5 f 0 ;  
         r a m _ c e l l [               9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 5 9 c 9 c a e ;  
         r a m _ c e l l [             1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 9 2 7 0 b 5 9 ;  
         r a m _ c e l l [             1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b c e 5 1 e c 9 ;  
         r a m _ c e l l [             1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 5 d 7 1 d a 6 ;  
         r a m _ c e l l [             1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 d 1 e 8 1 b 1 ;  
         r a m _ c e l l [             1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 d a 8 8 b 8 c ;  
         r a m _ c e l l [             1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 f e 3 a 9 7 d ;  
         r a m _ c e l l [             1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 e c f d 5 3 d ;  
         r a m _ c e l l [             1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 1 c 8 e 6 9 5 ;  
         r a m _ c e l l [             1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 d e d b b e 4 ;  
         r a m _ c e l l [             1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 f 0 a b c 6 a ;  
         r a m _ c e l l [             2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 1 1 4 6 c 5 0 ;  
         r a m _ c e l l [             2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 1 4 0 f 2 7 4 ;  
         r a m _ c e l l [             2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 8 c 0 1 6 6 6 ;  
         r a m _ c e l l [             2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 8 0 6 9 f 3 0 ;  
         r a m _ c e l l [             2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 7 1 5 1 a f b ;  
         r a m _ c e l l [             2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d a 8 3 e 7 a c ;  
         r a m _ c e l l [             2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 5 0 0 4 7 4 d ;  
         r a m _ c e l l [             2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 7 3 0 4 e 8 c ;  
         r a m _ c e l l [             2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f c 4 e 1 a 6 6 ;  
         r a m _ c e l l [             2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 3 6 c 2 d 6 6 ;  
         r a m _ c e l l [             3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 6 c d f 7 5 c ;  
         r a m _ c e l l [             3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 d 2 7 1 2 a c ;  
         r a m _ c e l l [             3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d d b f a 9 b b ;  
         r a m _ c e l l [             3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 8 2 5 5 c c 4 ;  
         r a m _ c e l l [             3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e b f 9 c 9 a 3 ;  
         r a m _ c e l l [             3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 1 7 2 5 1 e 5 ;  
         r a m _ c e l l [             3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 7 d 3 6 1 9 e ;  
         r a m _ c e l l [             3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 2 2 d b d 8 3 ;  
         r a m _ c e l l [             3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 3 2 1 a 2 0 a ;  
         r a m _ c e l l [             3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 4 0 9 0 e a a ;  
         r a m _ c e l l [             4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 6 8 b 0 3 7 9 ;  
         r a m _ c e l l [             4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 2 a 9 4 b 4 1 ;  
         r a m _ c e l l [             4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d a 0 3 4 4 3 d ;  
         r a m _ c e l l [             4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c b 3 e e 6 3 f ;  
         r a m _ c e l l [             4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 0 a 5 a b 9 f ;  
         r a m _ c e l l [             4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 b c 6 3 e 2 4 ;  
         r a m _ c e l l [             4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 2 9 5 c 6 d e ;  
         r a m _ c e l l [             4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 e c 7 5 9 3 0 ;  
         r a m _ c e l l [             4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d b 7 0 f 3 3 6 ;  
         r a m _ c e l l [             4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a c d 5 d d 7 c ;  
         r a m _ c e l l [             5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 2 d e 3 c a a ;  
         r a m _ c e l l [             5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 a f e b 3 4 e ;  
         r a m _ c e l l [             5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d b d e e a 5 9 ;  
         r a m _ c e l l [             5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 c 9 3 7 6 1 c ;  
         r a m _ c e l l [             5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 5 a f c 4 1 d ;  
         r a m _ c e l l [             5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 d b 6 a d 0 a ;  
         r a m _ c e l l [             5 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 5 5 d 1 0 8 c ;  
         r a m _ c e l l [             5 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 8 7 b 7 e 7 0 ;  
         r a m _ c e l l [             5 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 9 6 5 c 3 6 6 ;  
         r a m _ c e l l [             5 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 b 8 1 3 7 2 1 ;  
         r a m _ c e l l [             6 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f b 9 3 2 0 2 b ;  
         r a m _ c e l l [             6 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 7 9 7 2 0 7 4 ;  
         r a m _ c e l l [             6 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 3 c 7 b b c e ;  
         r a m _ c e l l [             6 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 7 6 2 8 1 0 e ;  
         / /   s r c   m a t r i x   A  
         r a m _ c e l l [             6 4 ]   =   3 2 ' h 9 0 6 5 6 7 a c ;  
         r a m _ c e l l [             6 5 ]   =   3 2 ' h 9 2 3 2 9 9 1 1 ;  
         r a m _ c e l l [             6 6 ]   =   3 2 ' h 8 2 7 6 c 2 e 1 ;  
         r a m _ c e l l [             6 7 ]   =   3 2 ' h a 3 4 c 8 6 d a ;  
         r a m _ c e l l [             6 8 ]   =   3 2 ' h 9 8 4 b 9 4 3 1 ;  
         r a m _ c e l l [             6 9 ]   =   3 2 ' h 3 c 6 f 8 0 d c ;  
         r a m _ c e l l [             7 0 ]   =   3 2 ' h b d b a d c 7 7 ;  
         r a m _ c e l l [             7 1 ]   =   3 2 ' h 3 5 7 c 0 6 a 6 ;  
         r a m _ c e l l [             7 2 ]   =   3 2 ' h c e 1 4 b e f c ;  
         r a m _ c e l l [             7 3 ]   =   3 2 ' h 5 f 1 8 b 4 b a ;  
         r a m _ c e l l [             7 4 ]   =   3 2 ' h 1 7 e 5 2 0 9 8 ;  
         r a m _ c e l l [             7 5 ]   =   3 2 ' h 7 3 b 7 f 6 d 4 ;  
         r a m _ c e l l [             7 6 ]   =   3 2 ' h 3 c e 3 b 8 c 6 ;  
         r a m _ c e l l [             7 7 ]   =   3 2 ' h 8 4 f 6 0 d c 9 ;  
         r a m _ c e l l [             7 8 ]   =   3 2 ' h 9 f a 7 0 3 8 8 ;  
         r a m _ c e l l [             7 9 ]   =   3 2 ' h c c a a 2 1 7 3 ;  
         r a m _ c e l l [             8 0 ]   =   3 2 ' h 7 5 0 8 f 8 4 f ;  
         r a m _ c e l l [             8 1 ]   =   3 2 ' h e e 0 6 e d 2 c ;  
         r a m _ c e l l [             8 2 ]   =   3 2 ' h c 6 0 4 3 2 2 a ;  
         r a m _ c e l l [             8 3 ]   =   3 2 ' h 7 8 b 5 d 5 5 c ;  
         r a m _ c e l l [             8 4 ]   =   3 2 ' h 0 0 a 2 1 7 8 c ;  
         r a m _ c e l l [             8 5 ]   =   3 2 ' h 7 9 b a 9 7 7 b ;  
         r a m _ c e l l [             8 6 ]   =   3 2 ' h 3 9 e 1 0 6 9 1 ;  
         r a m _ c e l l [             8 7 ]   =   3 2 ' h b 2 8 e a 2 4 d ;  
         r a m _ c e l l [             8 8 ]   =   3 2 ' h 0 f 3 4 2 d d 7 ;  
         r a m _ c e l l [             8 9 ]   =   3 2 ' h d d 3 e 2 8 1 6 ;  
         r a m _ c e l l [             9 0 ]   =   3 2 ' h 9 a d a 8 7 c 5 ;  
         r a m _ c e l l [             9 1 ]   =   3 2 ' h f 8 d 5 b 6 2 3 ;  
         r a m _ c e l l [             9 2 ]   =   3 2 ' h 2 4 8 2 5 a a d ;  
         r a m _ c e l l [             9 3 ]   =   3 2 ' h f d 3 b 8 a 2 2 ;  
         r a m _ c e l l [             9 4 ]   =   3 2 ' h a 3 9 d e b 8 2 ;  
         r a m _ c e l l [             9 5 ]   =   3 2 ' h f 6 9 b 1 5 b e ;  
         r a m _ c e l l [             9 6 ]   =   3 2 ' h e 7 f 8 4 f 8 7 ;  
         r a m _ c e l l [             9 7 ]   =   3 2 ' h f f 6 5 b 9 3 4 ;  
         r a m _ c e l l [             9 8 ]   =   3 2 ' h 2 4 7 4 b b a 2 ;  
         r a m _ c e l l [             9 9 ]   =   3 2 ' h 6 3 f 0 4 8 8 a ;  
         r a m _ c e l l [           1 0 0 ]   =   3 2 ' h 9 f 0 4 6 5 b 7 ;  
         r a m _ c e l l [           1 0 1 ]   =   3 2 ' h b a 0 8 f c 5 5 ;  
         r a m _ c e l l [           1 0 2 ]   =   3 2 ' h 3 7 6 d 9 a c a ;  
         r a m _ c e l l [           1 0 3 ]   =   3 2 ' h 7 9 f f 6 8 4 1 ;  
         r a m _ c e l l [           1 0 4 ]   =   3 2 ' h 4 b 8 7 9 b f 0 ;  
         r a m _ c e l l [           1 0 5 ]   =   3 2 ' h 6 1 b f d 7 d e ;  
         r a m _ c e l l [           1 0 6 ]   =   3 2 ' h 5 0 4 5 3 2 c d ;  
         r a m _ c e l l [           1 0 7 ]   =   3 2 ' h 1 3 2 a f e d 9 ;  
         r a m _ c e l l [           1 0 8 ]   =   3 2 ' h c 7 6 6 1 2 1 7 ;  
         r a m _ c e l l [           1 0 9 ]   =   3 2 ' h d f f d 2 2 a 1 ;  
         r a m _ c e l l [           1 1 0 ]   =   3 2 ' h b d a a 7 3 4 e ;  
         r a m _ c e l l [           1 1 1 ]   =   3 2 ' h 7 0 c b 6 3 e 6 ;  
         r a m _ c e l l [           1 1 2 ]   =   3 2 ' h 1 e 4 3 4 a 3 4 ;  
         r a m _ c e l l [           1 1 3 ]   =   3 2 ' h 5 a 5 b 7 d c 4 ;  
         r a m _ c e l l [           1 1 4 ]   =   3 2 ' h 5 0 a 9 4 6 d 4 ;  
         r a m _ c e l l [           1 1 5 ]   =   3 2 ' h f f 0 1 d 2 d 7 ;  
         r a m _ c e l l [           1 1 6 ]   =   3 2 ' h b d 2 5 d d f 7 ;  
         r a m _ c e l l [           1 1 7 ]   =   3 2 ' h f e 6 a 1 6 5 c ;  
         r a m _ c e l l [           1 1 8 ]   =   3 2 ' h f a 9 4 9 7 c a ;  
         r a m _ c e l l [           1 1 9 ]   =   3 2 ' h b 7 b 7 b 2 4 f ;  
         r a m _ c e l l [           1 2 0 ]   =   3 2 ' h 9 4 f 7 1 9 d f ;  
         r a m _ c e l l [           1 2 1 ]   =   3 2 ' h e 5 5 7 e f 3 5 ;  
         r a m _ c e l l [           1 2 2 ]   =   3 2 ' h 4 9 1 c 7 a 1 3 ;  
         r a m _ c e l l [           1 2 3 ]   =   3 2 ' h f 5 4 8 4 7 2 d ;  
         r a m _ c e l l [           1 2 4 ]   =   3 2 ' h c 0 4 5 6 4 8 f ;  
         r a m _ c e l l [           1 2 5 ]   =   3 2 ' h 3 4 c 0 c 3 7 e ;  
         r a m _ c e l l [           1 2 6 ]   =   3 2 ' h 2 4 b 6 1 5 f 6 ;  
         r a m _ c e l l [           1 2 7 ]   =   3 2 ' h 8 6 9 9 9 6 9 a ;  
         / /   s r c   m a t r i x   B  
         r a m _ c e l l [           1 2 8 ]   =   3 2 ' h d 8 6 e e 1 0 a ;  
         r a m _ c e l l [           1 2 9 ]   =   3 2 ' h a b c d b 2 b 6 ;  
         r a m _ c e l l [           1 3 0 ]   =   3 2 ' h a 7 4 9 3 0 f 0 ;  
         r a m _ c e l l [           1 3 1 ]   =   3 2 ' h 0 b 0 3 9 e d 8 ;  
         r a m _ c e l l [           1 3 2 ]   =   3 2 ' h 5 7 8 3 f 4 2 1 ;  
         r a m _ c e l l [           1 3 3 ]   =   3 2 ' h 2 b c b 9 c 5 5 ;  
         r a m _ c e l l [           1 3 4 ]   =   3 2 ' h 1 5 2 3 f 9 0 3 ;  
         r a m _ c e l l [           1 3 5 ]   =   3 2 ' h 5 f a 0 2 a 2 4 ;  
         r a m _ c e l l [           1 3 6 ]   =   3 2 ' h 5 c c 1 a 7 5 3 ;  
         r a m _ c e l l [           1 3 7 ]   =   3 2 ' h 2 b 6 7 9 1 e 2 ;  
         r a m _ c e l l [           1 3 8 ]   =   3 2 ' h 1 7 4 8 8 9 1 7 ;  
         r a m _ c e l l [           1 3 9 ]   =   3 2 ' h c e f 9 f 5 c b ;  
         r a m _ c e l l [           1 4 0 ]   =   3 2 ' h e d 0 c f b 5 1 ;  
         r a m _ c e l l [           1 4 1 ]   =   3 2 ' h 9 2 0 1 0 c 1 2 ;  
         r a m _ c e l l [           1 4 2 ]   =   3 2 ' h c e 5 7 3 f 8 2 ;  
         r a m _ c e l l [           1 4 3 ]   =   3 2 ' h e 9 3 f e 2 8 c ;  
         r a m _ c e l l [           1 4 4 ]   =   3 2 ' h f e 7 e e d 2 d ;  
         r a m _ c e l l [           1 4 5 ]   =   3 2 ' h 9 4 c 0 7 a e 1 ;  
         r a m _ c e l l [           1 4 6 ]   =   3 2 ' h 9 0 1 6 9 c 1 8 ;  
         r a m _ c e l l [           1 4 7 ]   =   3 2 ' h 7 f b a b 6 8 c ;  
         r a m _ c e l l [           1 4 8 ]   =   3 2 ' h e 6 b f 5 6 1 6 ;  
         r a m _ c e l l [           1 4 9 ]   =   3 2 ' h 3 2 8 e c 2 5 3 ;  
         r a m _ c e l l [           1 5 0 ]   =   3 2 ' h a 0 a 7 6 7 d b ;  
         r a m _ c e l l [           1 5 1 ]   =   3 2 ' h d 9 1 5 e 4 e 7 ;  
         r a m _ c e l l [           1 5 2 ]   =   3 2 ' h 7 9 4 5 9 2 9 5 ;  
         r a m _ c e l l [           1 5 3 ]   =   3 2 ' h 7 9 2 7 6 f 2 b ;  
         r a m _ c e l l [           1 5 4 ]   =   3 2 ' h e 9 c 9 4 c 9 7 ;  
         r a m _ c e l l [           1 5 5 ]   =   3 2 ' h 8 f 3 0 5 b 1 2 ;  
         r a m _ c e l l [           1 5 6 ]   =   3 2 ' h 1 7 2 d 6 2 3 a ;  
         r a m _ c e l l [           1 5 7 ]   =   3 2 ' h 7 9 0 2 1 c c 1 ;  
         r a m _ c e l l [           1 5 8 ]   =   3 2 ' h d c 8 7 2 b 2 7 ;  
         r a m _ c e l l [           1 5 9 ]   =   3 2 ' h 5 4 2 7 f 7 5 6 ;  
         r a m _ c e l l [           1 6 0 ]   =   3 2 ' h 6 c c 6 a b 4 3 ;  
         r a m _ c e l l [           1 6 1 ]   =   3 2 ' h c 4 7 c a f d 4 ;  
         r a m _ c e l l [           1 6 2 ]   =   3 2 ' h c c 5 c 5 4 f 0 ;  
         r a m _ c e l l [           1 6 3 ]   =   3 2 ' h f 3 a 9 3 3 9 c ;  
         r a m _ c e l l [           1 6 4 ]   =   3 2 ' h 9 7 2 4 6 d 6 5 ;  
         r a m _ c e l l [           1 6 5 ]   =   3 2 ' h f d e 2 e c 9 3 ;  
         r a m _ c e l l [           1 6 6 ]   =   3 2 ' h 5 e 6 c 3 b e d ;  
         r a m _ c e l l [           1 6 7 ]   =   3 2 ' h 7 b 1 a b d 6 3 ;  
         r a m _ c e l l [           1 6 8 ]   =   3 2 ' h 2 b b a 7 6 6 e ;  
         r a m _ c e l l [           1 6 9 ]   =   3 2 ' h 4 a 8 e b a b d ;  
         r a m _ c e l l [           1 7 0 ]   =   3 2 ' h 4 4 5 c 1 3 3 6 ;  
         r a m _ c e l l [           1 7 1 ]   =   3 2 ' h 4 c b 6 8 6 2 5 ;  
         r a m _ c e l l [           1 7 2 ]   =   3 2 ' h 0 d 4 1 3 d 5 c ;  
         r a m _ c e l l [           1 7 3 ]   =   3 2 ' h 0 7 7 0 d 1 d 1 ;  
         r a m _ c e l l [           1 7 4 ]   =   3 2 ' h 8 1 8 d 5 2 3 7 ;  
         r a m _ c e l l [           1 7 5 ]   =   3 2 ' h 6 9 1 6 4 c 1 0 ;  
         r a m _ c e l l [           1 7 6 ]   =   3 2 ' h c c 8 4 a 5 e 3 ;  
         r a m _ c e l l [           1 7 7 ]   =   3 2 ' h 9 5 e 1 0 c c f ;  
         r a m _ c e l l [           1 7 8 ]   =   3 2 ' h b e 4 b 4 7 b d ;  
         r a m _ c e l l [           1 7 9 ]   =   3 2 ' h 4 c 1 a f 3 1 f ;  
         r a m _ c e l l [           1 8 0 ]   =   3 2 ' h 6 4 5 3 5 4 f d ;  
         r a m _ c e l l [           1 8 1 ]   =   3 2 ' h 3 3 f d a a 1 8 ;  
         r a m _ c e l l [           1 8 2 ]   =   3 2 ' h 1 9 8 5 5 f d 9 ;  
         r a m _ c e l l [           1 8 3 ]   =   3 2 ' h 7 7 5 d 6 f d b ;  
         r a m _ c e l l [           1 8 4 ]   =   3 2 ' h 8 3 5 0 9 f 3 c ;  
         r a m _ c e l l [           1 8 5 ]   =   3 2 ' h f 0 2 9 e 1 0 b ;  
         r a m _ c e l l [           1 8 6 ]   =   3 2 ' h 8 f 4 7 8 8 6 3 ;  
         r a m _ c e l l [           1 8 7 ]   =   3 2 ' h 1 9 a 6 7 1 c 6 ;  
         r a m _ c e l l [           1 8 8 ]   =   3 2 ' h 6 c b 4 7 7 c a ;  
         r a m _ c e l l [           1 8 9 ]   =   3 2 ' h 9 8 f 1 f 0 3 c ;  
         r a m _ c e l l [           1 9 0 ]   =   3 2 ' h f 6 0 6 f e 2 5 ;  
         r a m _ c e l l [           1 9 1 ]   =   3 2 ' h c 8 c 1 8 e 3 b ;  
 e n d  
  
 e n d m o d u l e  
  
 