�� 
 m o d u l e   m e m   # (                                       / /    
         p a r a m e t e r     A D D R _ L E N     =   1 1       / /    
 )   (  
         i n p u t     c l k ,   r s t ,  
         i n p u t     [ A D D R _ L E N - 1 : 0 ]   a d d r ,   / /   m e m o r y   a d d r e s s  
         o u t p u t   r e g   [ 3 1 : 0 ]   r d _ d a t a ,     / /   d a t a   r e a d   o u t  
         i n p u t     w r _ r e q ,  
         i n p u t     [ 3 1 : 0 ]   w r _ d a t a               / /   d a t a   w r i t e   i n  
 ) ;  
 l o c a l p a r a m   M E M _ S I Z E   =   1 < < A D D R _ L E N ;  
 r e g   [ 3 1 : 0 ]   r a m _ c e l l   [ M E M _ S I Z E ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )  
                 r d _ d a t a   < =   0 ;  
         e l s e  
                 r d _ d a t a   < =   r a m _ c e l l [ a d d r ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k )  
         i f ( w r _ r e q )    
                 r a m _ c e l l [ a d d r ]   < =   w r _ d a t a ;  
  
 i n i t i a l   b e g i n  
         / /   d s t   m a t r i x   C  
         r a m _ c e l l [               0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 b 9 3 4 2 0 1 ;  
         r a m _ c e l l [               1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 6 6 2 a 3 d a ;  
         r a m _ c e l l [               2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 2 a 6 f e 4 0 ;  
         r a m _ c e l l [               3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 5 6 7 7 f b 2 ;  
         r a m _ c e l l [               4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 6 e 0 4 5 8 5 ;  
         r a m _ c e l l [               5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 9 a 2 f 2 b 8 ;  
         r a m _ c e l l [               6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 7 8 2 e 3 4 f ;  
         r a m _ c e l l [               7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 2 8 0 8 f c 8 ;  
         r a m _ c e l l [               8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 4 f 3 7 8 d a ;  
         r a m _ c e l l [               9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 5 f 6 2 9 7 4 ;  
         r a m _ c e l l [             1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 e b 2 2 e 5 2 ;  
         r a m _ c e l l [             1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 8 e d 9 1 d 9 ;  
         r a m _ c e l l [             1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 5 7 4 1 8 6 2 ;  
         r a m _ c e l l [             1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 2 1 8 6 0 e 1 ;  
         r a m _ c e l l [             1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 1 1 d 4 4 1 c ;  
         r a m _ c e l l [             1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 c a 0 4 6 0 3 ;  
         r a m _ c e l l [             1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 3 c b a c 0 9 ;  
         r a m _ c e l l [             1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 e 4 4 6 9 4 b ;  
         r a m _ c e l l [             1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 9 9 5 d 5 d 9 ;  
         r a m _ c e l l [             1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 5 2 e c 4 0 b ;  
         r a m _ c e l l [             2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 2 e 0 0 0 9 5 ;  
         r a m _ c e l l [             2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a f 2 4 c 3 9 0 ;  
         r a m _ c e l l [             2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 e 2 7 1 b b 0 ;  
         r a m _ c e l l [             2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 9 2 4 5 d 0 2 ;  
         r a m _ c e l l [             2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 4 d c d 4 7 e ;  
         r a m _ c e l l [             2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 6 3 1 c d 3 f ;  
         r a m _ c e l l [             2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e e 1 9 c a 5 9 ;  
         r a m _ c e l l [             2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 9 1 8 d 2 2 4 ;  
         r a m _ c e l l [             2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 e 6 4 4 a 8 0 ;  
         r a m _ c e l l [             2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 6 7 8 3 6 a 6 ;  
         r a m _ c e l l [             3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 1 6 7 a 2 2 d ;  
         r a m _ c e l l [             3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 a 6 9 7 8 f c ;  
         r a m _ c e l l [             3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 8 6 e 8 7 2 c ;  
         r a m _ c e l l [             3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 9 9 e d 2 4 f ;  
         r a m _ c e l l [             3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 a 6 0 1 3 c 9 ;  
         r a m _ c e l l [             3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 6 9 d 2 0 9 8 ;  
         r a m _ c e l l [             3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 9 4 8 9 1 9 5 ;  
         r a m _ c e l l [             3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 4 1 a c 3 9 d ;  
         r a m _ c e l l [             3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 4 8 2 c 5 1 a ;  
         r a m _ c e l l [             3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 2 6 d a 1 c d ;  
         r a m _ c e l l [             4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 6 c 2 d c 1 1 ;  
         r a m _ c e l l [             4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a a 0 c 1 2 f d ;  
         r a m _ c e l l [             4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 5 a e 4 7 e 8 ;  
         r a m _ c e l l [             4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 d f 3 4 9 3 b ;  
         r a m _ c e l l [             4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 6 b 0 7 7 c 2 ;  
         r a m _ c e l l [             4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e b 2 b 1 e 7 a ;  
         r a m _ c e l l [             4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 f 4 e c 4 7 1 ;  
         r a m _ c e l l [             4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 e a 2 4 0 b 0 ;  
         r a m _ c e l l [             4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 0 c 6 8 0 5 d ;  
         r a m _ c e l l [             4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 4 6 e 5 8 d 5 ;  
         r a m _ c e l l [             5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 5 2 0 f 4 0 b ;  
         r a m _ c e l l [             5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f f 5 6 b 0 5 5 ;  
         r a m _ c e l l [             5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 2 f c a f f f ;  
         r a m _ c e l l [             5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 7 8 1 0 8 e d ;  
         r a m _ c e l l [             5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 a 8 1 d c b 4 ;  
         r a m _ c e l l [             5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 c 3 8 c c 6 3 ;  
         r a m _ c e l l [             5 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 e 2 f 9 0 0 c ;  
         r a m _ c e l l [             5 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 8 1 b 0 5 8 3 ;  
         r a m _ c e l l [             5 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 c 5 d 2 a f b ;  
         r a m _ c e l l [             5 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 1 b 2 5 4 a b ;  
         r a m _ c e l l [             6 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 6 b f f f 6 8 ;  
         r a m _ c e l l [             6 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 1 d 9 7 f 4 2 ;  
         r a m _ c e l l [             6 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 e f 4 0 7 d 4 ;  
         r a m _ c e l l [             6 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 1 0 9 1 4 0 a ;  
         r a m _ c e l l [             6 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 4 7 4 f 5 c 5 ;  
         r a m _ c e l l [             6 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 6 4 9 3 0 c 1 ;  
         r a m _ c e l l [             6 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 e b 5 a 1 a 4 ;  
         r a m _ c e l l [             6 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 f b 1 2 e 4 f ;  
         r a m _ c e l l [             6 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 8 d 3 c e 0 4 ;  
         r a m _ c e l l [             6 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 1 2 e 3 c e 8 ;  
         r a m _ c e l l [             7 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 a 9 e 2 5 8 f ;  
         r a m _ c e l l [             7 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 4 d 4 9 f 1 0 ;  
         r a m _ c e l l [             7 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 e 6 a 0 d 9 1 ;  
         r a m _ c e l l [             7 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 9 3 8 2 8 1 2 ;  
         r a m _ c e l l [             7 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 2 1 9 8 5 7 1 ;  
         r a m _ c e l l [             7 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 7 8 f b 4 8 0 ;  
         r a m _ c e l l [             7 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 5 6 9 c b 0 1 ;  
         r a m _ c e l l [             7 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 6 4 a c 8 d c ;  
         r a m _ c e l l [             7 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 5 5 9 2 5 5 b ;  
         r a m _ c e l l [             7 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 4 5 2 2 b c b ;  
         r a m _ c e l l [             8 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 f 4 5 2 0 8 6 ;  
         r a m _ c e l l [             8 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 7 6 2 f 5 9 4 ;  
         r a m _ c e l l [             8 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 b 6 8 c 2 2 6 ;  
         r a m _ c e l l [             8 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 f 5 3 7 f b e ;  
         r a m _ c e l l [             8 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 1 1 1 6 a 2 0 ;  
         r a m _ c e l l [             8 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 9 f 3 9 0 d 7 ;  
         r a m _ c e l l [             8 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d f 6 c 6 2 e 3 ;  
         r a m _ c e l l [             8 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 8 d 9 6 a 0 9 ;  
         r a m _ c e l l [             8 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 7 f 5 9 4 d 6 ;  
         r a m _ c e l l [             8 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 c 1 4 3 9 0 a ;  
         r a m _ c e l l [             9 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 0 c d 0 b 0 4 ;  
         r a m _ c e l l [             9 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 f 3 8 8 c 9 c ;  
         r a m _ c e l l [             9 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 0 6 9 f 5 9 c ;  
         r a m _ c e l l [             9 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b a 2 4 6 a a c ;  
         r a m _ c e l l [             9 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 2 0 d 1 c 4 6 ;  
         r a m _ c e l l [             9 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 2 8 d 4 c 2 0 ;  
         r a m _ c e l l [             9 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 7 e 4 b 0 e d ;  
         r a m _ c e l l [             9 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a c a d 0 8 a 4 ;  
         r a m _ c e l l [             9 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 8 0 7 5 b 5 c ;  
         r a m _ c e l l [             9 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 6 f f d 4 a c ;  
         r a m _ c e l l [           1 0 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 7 e 8 b 7 5 5 ;  
         r a m _ c e l l [           1 0 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 6 6 2 1 a c 9 ;  
         r a m _ c e l l [           1 0 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 8 a 7 d d 6 9 ;  
         r a m _ c e l l [           1 0 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 8 f 1 4 2 6 6 ;  
         r a m _ c e l l [           1 0 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 4 a 5 7 9 f c ;  
         r a m _ c e l l [           1 0 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 2 2 6 9 9 a 5 ;  
         r a m _ c e l l [           1 0 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 d 4 0 5 8 4 3 ;  
         r a m _ c e l l [           1 0 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 2 c 0 d 5 9 5 ;  
         r a m _ c e l l [           1 0 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 d 6 9 1 e 7 0 ;  
         r a m _ c e l l [           1 0 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 f 2 d 7 b f e ;  
         r a m _ c e l l [           1 1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d a 7 9 b 7 e d ;  
         r a m _ c e l l [           1 1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c a 2 7 5 0 e 7 ;  
         r a m _ c e l l [           1 1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 c 2 0 1 7 2 0 ;  
         r a m _ c e l l [           1 1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 5 b f 7 6 0 8 ;  
         r a m _ c e l l [           1 1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 d d 7 4 b a 8 ;  
         r a m _ c e l l [           1 1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 3 f 7 e 5 0 6 ;  
         r a m _ c e l l [           1 1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 5 0 3 2 a 6 b ;  
         r a m _ c e l l [           1 1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 2 c 5 a 6 8 b ;  
         r a m _ c e l l [           1 1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 4 6 2 c 0 7 8 ;  
         r a m _ c e l l [           1 1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 5 1 8 3 e 5 9 ;  
         r a m _ c e l l [           1 2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 9 0 d 5 b 9 f ;  
         r a m _ c e l l [           1 2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 5 4 8 2 6 a f ;  
         r a m _ c e l l [           1 2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 f 7 4 7 c 9 e ;  
         r a m _ c e l l [           1 2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 e 9 9 3 4 7 e ;  
         r a m _ c e l l [           1 2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 c 8 8 e 6 1 4 ;  
         r a m _ c e l l [           1 2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 6 e b 1 c 3 4 ;  
         r a m _ c e l l [           1 2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 3 8 1 1 d b 3 ;  
         r a m _ c e l l [           1 2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 3 b 4 9 0 0 8 ;  
         r a m _ c e l l [           1 2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 e 2 3 7 0 d b ;  
         r a m _ c e l l [           1 2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 c a 9 2 5 4 3 ;  
         r a m _ c e l l [           1 3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 e 7 c 3 2 6 7 ;  
         r a m _ c e l l [           1 3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 f a 5 6 3 7 f ;  
         r a m _ c e l l [           1 3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 3 d 3 2 3 c 9 ;  
         r a m _ c e l l [           1 3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 8 2 1 e 6 a 1 ;  
         r a m _ c e l l [           1 3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 d 3 e 7 4 f 4 ;  
         r a m _ c e l l [           1 3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c d e 1 f f 3 c ;  
         r a m _ c e l l [           1 3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 1 1 5 b 1 d 9 ;  
         r a m _ c e l l [           1 3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 7 8 5 f e 6 b ;  
         r a m _ c e l l [           1 3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 9 2 9 2 2 5 7 ;  
         r a m _ c e l l [           1 3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 7 2 5 a e a 9 ;  
         r a m _ c e l l [           1 4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 7 5 9 8 9 9 0 ;  
         r a m _ c e l l [           1 4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 4 8 b b 6 8 7 ;  
         r a m _ c e l l [           1 4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 2 3 9 2 5 2 d ;  
         r a m _ c e l l [           1 4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 4 c d 8 8 1 f ;  
         r a m _ c e l l [           1 4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 8 2 f 1 9 3 4 ;  
         r a m _ c e l l [           1 4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 a 8 b 0 0 f f ;  
         r a m _ c e l l [           1 4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 1 3 f 7 6 3 3 ;  
         r a m _ c e l l [           1 4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 c d 9 f d c 8 ;  
         r a m _ c e l l [           1 4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 0 1 4 d 6 3 d ;  
         r a m _ c e l l [           1 4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 9 c 1 4 a 0 6 ;  
         r a m _ c e l l [           1 5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 d e 2 4 5 3 2 ;  
         r a m _ c e l l [           1 5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 1 c 5 8 3 c d ;  
         r a m _ c e l l [           1 5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 4 7 a 6 3 9 c ;  
         r a m _ c e l l [           1 5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 0 0 6 8 2 4 3 ;  
         r a m _ c e l l [           1 5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 7 9 2 e 6 5 3 ;  
         r a m _ c e l l [           1 5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 c d 3 5 f 8 b ;  
         r a m _ c e l l [           1 5 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 9 4 9 4 b 8 3 ;  
         r a m _ c e l l [           1 5 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 2 9 1 4 0 b 8 ;  
         r a m _ c e l l [           1 5 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 5 9 0 0 e d 8 ;  
         r a m _ c e l l [           1 5 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 4 7 2 4 f d 8 ;  
         r a m _ c e l l [           1 6 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 3 a f 7 9 4 1 ;  
         r a m _ c e l l [           1 6 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 0 d 7 8 0 d c ;  
         r a m _ c e l l [           1 6 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 5 d 4 3 a 5 e ;  
         r a m _ c e l l [           1 6 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 2 2 c 5 4 1 2 ;  
         r a m _ c e l l [           1 6 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 a 0 2 f 3 c b ;  
         r a m _ c e l l [           1 6 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 f 4 a 0 6 3 e ;  
         r a m _ c e l l [           1 6 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 e 0 7 1 5 f 8 ;  
         r a m _ c e l l [           1 6 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c d b 4 f 4 c 1 ;  
         r a m _ c e l l [           1 6 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 8 e 7 7 d 7 c ;  
         r a m _ c e l l [           1 6 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 0 3 b 0 6 1 5 ;  
         r a m _ c e l l [           1 7 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 e 8 1 a b 6 a ;  
         r a m _ c e l l [           1 7 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 6 4 b 5 b 1 4 ;  
         r a m _ c e l l [           1 7 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 a a 1 0 8 1 7 ;  
         r a m _ c e l l [           1 7 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 5 f f 5 2 d 8 ;  
         r a m _ c e l l [           1 7 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 4 1 3 c 1 8 c ;  
         r a m _ c e l l [           1 7 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 2 6 f e c f e ;  
         r a m _ c e l l [           1 7 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 8 b 7 5 2 f 1 ;  
         r a m _ c e l l [           1 7 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 7 e 3 c d 8 4 ;  
         r a m _ c e l l [           1 7 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 6 d 5 b 5 2 a ;  
         r a m _ c e l l [           1 7 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 c a b a a 3 0 ;  
         r a m _ c e l l [           1 8 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 6 1 3 2 e f 1 ;  
         r a m _ c e l l [           1 8 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 f e c 7 1 d e ;  
         r a m _ c e l l [           1 8 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 0 9 a 6 8 5 6 ;  
         r a m _ c e l l [           1 8 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 2 1 5 2 0 2 a ;  
         r a m _ c e l l [           1 8 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 a 2 b 3 b 8 6 ;  
         r a m _ c e l l [           1 8 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 3 a 2 8 a 5 7 ;  
         r a m _ c e l l [           1 8 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 4 6 e f 4 5 4 ;  
         r a m _ c e l l [           1 8 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 1 6 9 b 7 7 1 ;  
         r a m _ c e l l [           1 8 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 2 a e 2 6 e c ;  
         r a m _ c e l l [           1 8 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e e 0 2 4 0 f 0 ;  
         r a m _ c e l l [           1 9 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 0 0 2 3 0 6 0 ;  
         r a m _ c e l l [           1 9 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c f 6 d 8 7 8 5 ;  
         r a m _ c e l l [           1 9 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 3 c d 5 1 a 4 ;  
         r a m _ c e l l [           1 9 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 9 6 6 c 5 1 a ;  
         r a m _ c e l l [           1 9 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 9 d f c f 5 8 ;  
         r a m _ c e l l [           1 9 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 1 5 2 f e 4 4 ;  
         r a m _ c e l l [           1 9 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 5 5 e d 3 6 9 ;  
         r a m _ c e l l [           1 9 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e a 7 3 b 9 b 1 ;  
         r a m _ c e l l [           1 9 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 2 d 7 d 7 3 4 ;  
         r a m _ c e l l [           1 9 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 c d 8 2 b f 6 ;  
         r a m _ c e l l [           2 0 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a e 5 5 7 9 0 7 ;  
         r a m _ c e l l [           2 0 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 5 f a 0 2 7 3 ;  
         r a m _ c e l l [           2 0 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 1 2 2 b 7 5 9 ;  
         r a m _ c e l l [           2 0 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 2 d 5 2 f f 5 ;  
         r a m _ c e l l [           2 0 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 d c 0 0 3 a f ;  
         r a m _ c e l l [           2 0 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 f a 8 2 9 4 5 ;  
         r a m _ c e l l [           2 0 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b b f a c 5 4 0 ;  
         r a m _ c e l l [           2 0 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 1 2 0 a e 2 e ;  
         r a m _ c e l l [           2 0 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 0 9 5 6 d c 8 ;  
         r a m _ c e l l [           2 0 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 5 0 e 1 e 2 c ;  
         r a m _ c e l l [           2 1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 6 8 e e c c 8 ;  
         r a m _ c e l l [           2 1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 9 1 f 1 7 c 7 ;  
         r a m _ c e l l [           2 1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a c 2 4 6 a 5 1 ;  
         r a m _ c e l l [           2 1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 d 4 9 1 1 4 3 ;  
         r a m _ c e l l [           2 1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e c 0 d a c 1 d ;  
         r a m _ c e l l [           2 1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 7 3 b 2 b 1 e ;  
         r a m _ c e l l [           2 1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 f 2 e 1 0 4 c ;  
         r a m _ c e l l [           2 1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 6 f 6 c 4 5 9 ;  
         r a m _ c e l l [           2 1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 1 7 4 9 9 a 7 ;  
         r a m _ c e l l [           2 1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 1 d 0 e 8 2 4 ;  
         r a m _ c e l l [           2 2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 f 0 7 5 a 2 f ;  
         r a m _ c e l l [           2 2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 6 3 c 6 9 4 5 ;  
         r a m _ c e l l [           2 2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 a e 7 d 6 2 8 ;  
         r a m _ c e l l [           2 2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 1 b b a 9 a 6 ;  
         r a m _ c e l l [           2 2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 5 f 0 f 6 6 2 ;  
         r a m _ c e l l [           2 2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 6 5 f f e 7 5 ;  
         r a m _ c e l l [           2 2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 4 8 9 5 e c 0 ;  
         r a m _ c e l l [           2 2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 6 0 6 f a d 3 ;  
         r a m _ c e l l [           2 2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 7 f 3 9 c d b ;  
         r a m _ c e l l [           2 2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 e 4 1 f b 1 2 ;  
         r a m _ c e l l [           2 3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 b d e 5 3 c d ;  
         r a m _ c e l l [           2 3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 8 0 4 c 3 f 0 ;  
         r a m _ c e l l [           2 3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 7 0 9 c d 3 c ;  
         r a m _ c e l l [           2 3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 3 e b 3 6 7 c ;  
         r a m _ c e l l [           2 3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b d 6 9 5 2 f 5 ;  
         r a m _ c e l l [           2 3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 f 5 1 3 2 2 1 ;  
         r a m _ c e l l [           2 3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 5 f 5 c 3 2 d ;  
         r a m _ c e l l [           2 3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f e 7 3 d 9 d e ;  
         r a m _ c e l l [           2 3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 2 2 8 e a 0 6 ;  
         r a m _ c e l l [           2 3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 6 4 2 8 e f 1 ;  
         r a m _ c e l l [           2 4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 e 4 3 0 d f f ;  
         r a m _ c e l l [           2 4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 1 4 b 9 5 c 5 ;  
         r a m _ c e l l [           2 4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 5 4 3 8 e d f ;  
         r a m _ c e l l [           2 4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 f 5 4 b 5 b c ;  
         r a m _ c e l l [           2 4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 1 e 9 4 f 7 5 ;  
         r a m _ c e l l [           2 4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 3 0 8 1 c 7 3 ;  
         r a m _ c e l l [           2 4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 f 3 6 4 b 8 9 ;  
         r a m _ c e l l [           2 4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 a a 7 e 9 1 2 ;  
         r a m _ c e l l [           2 4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 f 9 1 9 9 7 f ;  
         r a m _ c e l l [           2 4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 5 6 9 f f 7 4 ;  
         r a m _ c e l l [           2 5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 1 9 c d 8 0 8 ;  
         r a m _ c e l l [           2 5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 9 e e a 3 f a ;  
         r a m _ c e l l [           2 5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 5 6 3 e 4 f e ;  
         r a m _ c e l l [           2 5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 0 0 6 c f 6 1 ;  
         r a m _ c e l l [           2 5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 9 a b 7 c 9 d ;  
         r a m _ c e l l [           2 5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 0 b 1 1 c 3 a ;  
         / /   s r c   m a t r i x   A  
         r a m _ c e l l [           2 5 6 ]   =   3 2 ' h 1 1 2 d b f 5 3 ;  
         r a m _ c e l l [           2 5 7 ]   =   3 2 ' h f c a 8 9 b 6 b ;  
         r a m _ c e l l [           2 5 8 ]   =   3 2 ' h 8 7 d 1 8 2 1 e ;  
         r a m _ c e l l [           2 5 9 ]   =   3 2 ' h 1 9 b 9 6 8 2 3 ;  
         r a m _ c e l l [           2 6 0 ]   =   3 2 ' h 3 b c 1 4 b f c ;  
         r a m _ c e l l [           2 6 1 ]   =   3 2 ' h d f 2 e f 4 d 7 ;  
         r a m _ c e l l [           2 6 2 ]   =   3 2 ' h 3 c 0 4 1 3 f 0 ;  
         r a m _ c e l l [           2 6 3 ]   =   3 2 ' h 4 c c 5 6 a 1 0 ;  
         r a m _ c e l l [           2 6 4 ]   =   3 2 ' h c a a e 7 e 9 7 ;  
         r a m _ c e l l [           2 6 5 ]   =   3 2 ' h 7 6 6 b a 9 6 1 ;  
         r a m _ c e l l [           2 6 6 ]   =   3 2 ' h c f 5 d 8 4 9 9 ;  
         r a m _ c e l l [           2 6 7 ]   =   3 2 ' h 0 4 b 4 8 4 d c ;  
         r a m _ c e l l [           2 6 8 ]   =   3 2 ' h e 9 a 4 e 2 b b ;  
         r a m _ c e l l [           2 6 9 ]   =   3 2 ' h 7 d b 9 7 0 2 7 ;  
         r a m _ c e l l [           2 7 0 ]   =   3 2 ' h 7 2 5 3 6 6 6 a ;  
         r a m _ c e l l [           2 7 1 ]   =   3 2 ' h 6 5 a d 5 2 c d ;  
         r a m _ c e l l [           2 7 2 ]   =   3 2 ' h 6 1 d c 5 7 3 a ;  
         r a m _ c e l l [           2 7 3 ]   =   3 2 ' h f 9 6 d a 0 3 e ;  
         r a m _ c e l l [           2 7 4 ]   =   3 2 ' h 3 a 9 0 7 c 9 a ;  
         r a m _ c e l l [           2 7 5 ]   =   3 2 ' h 6 8 1 8 d d 9 a ;  
         r a m _ c e l l [           2 7 6 ]   =   3 2 ' h 2 f b 1 6 a 2 7 ;  
         r a m _ c e l l [           2 7 7 ]   =   3 2 ' h f 5 8 9 5 2 4 a ;  
         r a m _ c e l l [           2 7 8 ]   =   3 2 ' h 3 0 5 a 0 c 8 0 ;  
         r a m _ c e l l [           2 7 9 ]   =   3 2 ' h 8 4 4 5 8 a c 0 ;  
         r a m _ c e l l [           2 8 0 ]   =   3 2 ' h 7 1 0 0 5 5 4 7 ;  
         r a m _ c e l l [           2 8 1 ]   =   3 2 ' h 5 f 1 1 0 e 7 f ;  
         r a m _ c e l l [           2 8 2 ]   =   3 2 ' h 8 0 b d 0 c f 2 ;  
         r a m _ c e l l [           2 8 3 ]   =   3 2 ' h f 9 1 a 3 6 8 c ;  
         r a m _ c e l l [           2 8 4 ]   =   3 2 ' h 4 3 4 6 e 5 3 b ;  
         r a m _ c e l l [           2 8 5 ]   =   3 2 ' h 8 1 3 9 1 3 9 2 ;  
         r a m _ c e l l [           2 8 6 ]   =   3 2 ' h b f 7 7 9 8 0 4 ;  
         r a m _ c e l l [           2 8 7 ]   =   3 2 ' h c f f 6 e 2 8 f ;  
         r a m _ c e l l [           2 8 8 ]   =   3 2 ' h 1 0 a 6 0 9 2 4 ;  
         r a m _ c e l l [           2 8 9 ]   =   3 2 ' h 3 0 3 e 0 0 f f ;  
         r a m _ c e l l [           2 9 0 ]   =   3 2 ' h 8 9 1 d d d 4 9 ;  
         r a m _ c e l l [           2 9 1 ]   =   3 2 ' h c b 2 4 c 1 0 f ;  
         r a m _ c e l l [           2 9 2 ]   =   3 2 ' h 7 6 c 6 e a 1 4 ;  
         r a m _ c e l l [           2 9 3 ]   =   3 2 ' h 8 e d 2 a a 8 7 ;  
         r a m _ c e l l [           2 9 4 ]   =   3 2 ' h 7 e b e e c 6 a ;  
         r a m _ c e l l [           2 9 5 ]   =   3 2 ' h d 3 c f 0 7 b 3 ;  
         r a m _ c e l l [           2 9 6 ]   =   3 2 ' h 7 0 0 1 7 1 5 7 ;  
         r a m _ c e l l [           2 9 7 ]   =   3 2 ' h e 2 9 1 9 d 1 5 ;  
         r a m _ c e l l [           2 9 8 ]   =   3 2 ' h 5 0 a a 2 6 8 f ;  
         r a m _ c e l l [           2 9 9 ]   =   3 2 ' h 3 b 2 8 7 4 8 0 ;  
         r a m _ c e l l [           3 0 0 ]   =   3 2 ' h 2 d f a 4 7 3 5 ;  
         r a m _ c e l l [           3 0 1 ]   =   3 2 ' h d 1 c 5 6 5 4 6 ;  
         r a m _ c e l l [           3 0 2 ]   =   3 2 ' h b 4 2 e d b 4 7 ;  
         r a m _ c e l l [           3 0 3 ]   =   3 2 ' h 7 9 6 c 7 1 1 9 ;  
         r a m _ c e l l [           3 0 4 ]   =   3 2 ' h 3 a f 9 7 3 4 1 ;  
         r a m _ c e l l [           3 0 5 ]   =   3 2 ' h 0 7 9 7 4 6 a a ;  
         r a m _ c e l l [           3 0 6 ]   =   3 2 ' h 2 3 8 4 d 3 1 9 ;  
         r a m _ c e l l [           3 0 7 ]   =   3 2 ' h 0 0 4 3 e 0 b 7 ;  
         r a m _ c e l l [           3 0 8 ]   =   3 2 ' h b b f 5 a b 8 8 ;  
         r a m _ c e l l [           3 0 9 ]   =   3 2 ' h d f c b 7 3 a 6 ;  
         r a m _ c e l l [           3 1 0 ]   =   3 2 ' h a 1 f 4 0 5 5 f ;  
         r a m _ c e l l [           3 1 1 ]   =   3 2 ' h b 6 e 2 3 f e 1 ;  
         r a m _ c e l l [           3 1 2 ]   =   3 2 ' h c 4 8 c 3 d 8 6 ;  
         r a m _ c e l l [           3 1 3 ]   =   3 2 ' h 2 0 9 0 6 1 b e ;  
         r a m _ c e l l [           3 1 4 ]   =   3 2 ' h e 8 e 0 2 c 4 8 ;  
         r a m _ c e l l [           3 1 5 ]   =   3 2 ' h 6 0 5 b 0 4 7 8 ;  
         r a m _ c e l l [           3 1 6 ]   =   3 2 ' h f a 2 c 2 a 8 b ;  
         r a m _ c e l l [           3 1 7 ]   =   3 2 ' h 2 2 e 6 3 8 e e ;  
         r a m _ c e l l [           3 1 8 ]   =   3 2 ' h 0 1 0 c 6 b 3 1 ;  
         r a m _ c e l l [           3 1 9 ]   =   3 2 ' h 1 7 e b 5 4 f b ;  
         r a m _ c e l l [           3 2 0 ]   =   3 2 ' h 9 3 2 c 0 2 8 8 ;  
         r a m _ c e l l [           3 2 1 ]   =   3 2 ' h 4 2 a 2 9 d 4 5 ;  
         r a m _ c e l l [           3 2 2 ]   =   3 2 ' h 9 a 6 5 5 f 7 9 ;  
         r a m _ c e l l [           3 2 3 ]   =   3 2 ' h b a a 8 9 b e 5 ;  
         r a m _ c e l l [           3 2 4 ]   =   3 2 ' h 2 1 6 c f 9 1 8 ;  
         r a m _ c e l l [           3 2 5 ]   =   3 2 ' h f 1 a b 6 6 1 7 ;  
         r a m _ c e l l [           3 2 6 ]   =   3 2 ' h 1 e 6 0 f 5 a 8 ;  
         r a m _ c e l l [           3 2 7 ]   =   3 2 ' h b e b a 2 b 0 0 ;  
         r a m _ c e l l [           3 2 8 ]   =   3 2 ' h 3 7 c 6 e 8 d 7 ;  
         r a m _ c e l l [           3 2 9 ]   =   3 2 ' h 7 e 1 f 6 0 d 1 ;  
         r a m _ c e l l [           3 3 0 ]   =   3 2 ' h f 3 d c 6 2 1 f ;  
         r a m _ c e l l [           3 3 1 ]   =   3 2 ' h 8 b f 3 a d c d ;  
         r a m _ c e l l [           3 3 2 ]   =   3 2 ' h 0 7 c 0 5 7 c 8 ;  
         r a m _ c e l l [           3 3 3 ]   =   3 2 ' h 8 7 4 0 9 8 5 f ;  
         r a m _ c e l l [           3 3 4 ]   =   3 2 ' h d 4 4 7 1 0 f d ;  
         r a m _ c e l l [           3 3 5 ]   =   3 2 ' h 3 4 3 3 d e 3 f ;  
         r a m _ c e l l [           3 3 6 ]   =   3 2 ' h 8 7 f b f 9 b 6 ;  
         r a m _ c e l l [           3 3 7 ]   =   3 2 ' h a 8 0 a 2 0 4 e ;  
         r a m _ c e l l [           3 3 8 ]   =   3 2 ' h b 2 6 6 9 e f 0 ;  
         r a m _ c e l l [           3 3 9 ]   =   3 2 ' h 9 c 6 2 7 7 9 c ;  
         r a m _ c e l l [           3 4 0 ]   =   3 2 ' h d b 0 5 8 c 8 a ;  
         r a m _ c e l l [           3 4 1 ]   =   3 2 ' h 3 b 5 2 5 b 8 a ;  
         r a m _ c e l l [           3 4 2 ]   =   3 2 ' h d 8 4 f 4 b a a ;  
         r a m _ c e l l [           3 4 3 ]   =   3 2 ' h a d 5 d 6 4 c e ;  
         r a m _ c e l l [           3 4 4 ]   =   3 2 ' h c 0 2 0 a 1 1 6 ;  
         r a m _ c e l l [           3 4 5 ]   =   3 2 ' h 3 1 8 c d 4 4 d ;  
         r a m _ c e l l [           3 4 6 ]   =   3 2 ' h 3 7 8 3 6 1 c 2 ;  
         r a m _ c e l l [           3 4 7 ]   =   3 2 ' h 4 9 6 0 e a 6 e ;  
         r a m _ c e l l [           3 4 8 ]   =   3 2 ' h 8 a b f 5 5 9 9 ;  
         r a m _ c e l l [           3 4 9 ]   =   3 2 ' h 4 b c 1 f 6 c 9 ;  
         r a m _ c e l l [           3 5 0 ]   =   3 2 ' h 1 a c 3 7 d e b ;  
         r a m _ c e l l [           3 5 1 ]   =   3 2 ' h f 9 b a c 4 6 0 ;  
         r a m _ c e l l [           3 5 2 ]   =   3 2 ' h e d f e d 9 9 9 ;  
         r a m _ c e l l [           3 5 3 ]   =   3 2 ' h 4 7 f a 8 8 7 a ;  
         r a m _ c e l l [           3 5 4 ]   =   3 2 ' h d 8 a b 1 9 a 4 ;  
         r a m _ c e l l [           3 5 5 ]   =   3 2 ' h 7 f 7 4 6 5 4 b ;  
         r a m _ c e l l [           3 5 6 ]   =   3 2 ' h 3 6 d 1 f 2 8 8 ;  
         r a m _ c e l l [           3 5 7 ]   =   3 2 ' h 3 2 4 f 0 7 d d ;  
         r a m _ c e l l [           3 5 8 ]   =   3 2 ' h 5 e 2 9 c 4 0 1 ;  
         r a m _ c e l l [           3 5 9 ]   =   3 2 ' h 0 0 3 a a 4 7 0 ;  
         r a m _ c e l l [           3 6 0 ]   =   3 2 ' h 2 b 6 9 b 7 6 5 ;  
         r a m _ c e l l [           3 6 1 ]   =   3 2 ' h 3 5 0 f e e f 0 ;  
         r a m _ c e l l [           3 6 2 ]   =   3 2 ' h e 1 9 7 f 6 c 2 ;  
         r a m _ c e l l [           3 6 3 ]   =   3 2 ' h e c 6 e 9 2 b 6 ;  
         r a m _ c e l l [           3 6 4 ]   =   3 2 ' h a 0 a 9 4 8 f c ;  
         r a m _ c e l l [           3 6 5 ]   =   3 2 ' h 9 8 7 0 a 5 4 9 ;  
         r a m _ c e l l [           3 6 6 ]   =   3 2 ' h 6 c 7 1 9 4 c b ;  
         r a m _ c e l l [           3 6 7 ]   =   3 2 ' h 9 b b 9 e 4 b 1 ;  
         r a m _ c e l l [           3 6 8 ]   =   3 2 ' h b 1 6 f 6 c 3 0 ;  
         r a m _ c e l l [           3 6 9 ]   =   3 2 ' h 7 e 5 9 3 b 8 4 ;  
         r a m _ c e l l [           3 7 0 ]   =   3 2 ' h 7 1 d 9 2 c 9 3 ;  
         r a m _ c e l l [           3 7 1 ]   =   3 2 ' h b 7 2 7 0 c 4 5 ;  
         r a m _ c e l l [           3 7 2 ]   =   3 2 ' h 5 5 7 a b 4 4 1 ;  
         r a m _ c e l l [           3 7 3 ]   =   3 2 ' h 7 a d c 9 f f 3 ;  
         r a m _ c e l l [           3 7 4 ]   =   3 2 ' h d 2 5 7 2 c 8 2 ;  
         r a m _ c e l l [           3 7 5 ]   =   3 2 ' h e c 5 3 3 b f e ;  
         r a m _ c e l l [           3 7 6 ]   =   3 2 ' h 7 a a 4 e d c 4 ;  
         r a m _ c e l l [           3 7 7 ]   =   3 2 ' h f b 0 3 e 0 4 4 ;  
         r a m _ c e l l [           3 7 8 ]   =   3 2 ' h 7 7 c 4 0 6 9 e ;  
         r a m _ c e l l [           3 7 9 ]   =   3 2 ' h 2 0 d 1 3 6 1 2 ;  
         r a m _ c e l l [           3 8 0 ]   =   3 2 ' h a 4 c d e 8 7 c ;  
         r a m _ c e l l [           3 8 1 ]   =   3 2 ' h a a 5 f 3 d 2 0 ;  
         r a m _ c e l l [           3 8 2 ]   =   3 2 ' h 0 7 9 a 3 b 9 b ;  
         r a m _ c e l l [           3 8 3 ]   =   3 2 ' h 5 6 4 8 5 2 2 7 ;  
         r a m _ c e l l [           3 8 4 ]   =   3 2 ' h 2 0 9 7 6 3 1 9 ;  
         r a m _ c e l l [           3 8 5 ]   =   3 2 ' h 0 1 8 5 6 2 0 3 ;  
         r a m _ c e l l [           3 8 6 ]   =   3 2 ' h b b 3 e 2 f 7 3 ;  
         r a m _ c e l l [           3 8 7 ]   =   3 2 ' h a 2 7 e a e 8 d ;  
         r a m _ c e l l [           3 8 8 ]   =   3 2 ' h c 3 4 a 2 6 c 6 ;  
         r a m _ c e l l [           3 8 9 ]   =   3 2 ' h 4 a 7 e 1 0 a b ;  
         r a m _ c e l l [           3 9 0 ]   =   3 2 ' h 3 e 7 0 7 c b 6 ;  
         r a m _ c e l l [           3 9 1 ]   =   3 2 ' h 1 6 b b 6 5 f c ;  
         r a m _ c e l l [           3 9 2 ]   =   3 2 ' h f 4 4 0 2 f 5 0 ;  
         r a m _ c e l l [           3 9 3 ]   =   3 2 ' h 4 f 5 0 e 1 1 9 ;  
         r a m _ c e l l [           3 9 4 ]   =   3 2 ' h 1 9 1 8 5 3 3 2 ;  
         r a m _ c e l l [           3 9 5 ]   =   3 2 ' h a f f 1 9 4 4 b ;  
         r a m _ c e l l [           3 9 6 ]   =   3 2 ' h c f b a a b 3 1 ;  
         r a m _ c e l l [           3 9 7 ]   =   3 2 ' h a 7 f 0 5 0 0 b ;  
         r a m _ c e l l [           3 9 8 ]   =   3 2 ' h 2 0 d 2 7 2 b e ;  
         r a m _ c e l l [           3 9 9 ]   =   3 2 ' h d c d 1 5 2 3 e ;  
         r a m _ c e l l [           4 0 0 ]   =   3 2 ' h e f 1 c c 2 1 1 ;  
         r a m _ c e l l [           4 0 1 ]   =   3 2 ' h b 7 a 9 4 0 c b ;  
         r a m _ c e l l [           4 0 2 ]   =   3 2 ' h 8 6 c 4 7 9 6 4 ;  
         r a m _ c e l l [           4 0 3 ]   =   3 2 ' h 9 9 1 8 3 0 8 e ;  
         r a m _ c e l l [           4 0 4 ]   =   3 2 ' h c 3 a 8 b 6 6 2 ;  
         r a m _ c e l l [           4 0 5 ]   =   3 2 ' h 4 1 7 a 3 f 8 4 ;  
         r a m _ c e l l [           4 0 6 ]   =   3 2 ' h c 3 b d e a 6 9 ;  
         r a m _ c e l l [           4 0 7 ]   =   3 2 ' h 2 1 1 1 6 8 3 c ;  
         r a m _ c e l l [           4 0 8 ]   =   3 2 ' h 8 e 5 1 6 c 5 c ;  
         r a m _ c e l l [           4 0 9 ]   =   3 2 ' h c e f 3 9 3 b e ;  
         r a m _ c e l l [           4 1 0 ]   =   3 2 ' h 6 0 0 b 9 1 5 3 ;  
         r a m _ c e l l [           4 1 1 ]   =   3 2 ' h f d 0 f c 7 a e ;  
         r a m _ c e l l [           4 1 2 ]   =   3 2 ' h 7 2 e d c f 2 7 ;  
         r a m _ c e l l [           4 1 3 ]   =   3 2 ' h 1 3 9 2 3 9 e 0 ;  
         r a m _ c e l l [           4 1 4 ]   =   3 2 ' h 1 3 9 b 1 4 e 4 ;  
         r a m _ c e l l [           4 1 5 ]   =   3 2 ' h 1 7 6 e f 5 6 6 ;  
         r a m _ c e l l [           4 1 6 ]   =   3 2 ' h 3 a 5 6 7 b c b ;  
         r a m _ c e l l [           4 1 7 ]   =   3 2 ' h 9 e 8 b 0 0 f f ;  
         r a m _ c e l l [           4 1 8 ]   =   3 2 ' h 4 4 9 8 a 3 7 8 ;  
         r a m _ c e l l [           4 1 9 ]   =   3 2 ' h 4 8 a 5 8 e 6 b ;  
         r a m _ c e l l [           4 2 0 ]   =   3 2 ' h a 0 8 7 b 8 1 e ;  
         r a m _ c e l l [           4 2 1 ]   =   3 2 ' h f f 1 6 8 f 7 2 ;  
         r a m _ c e l l [           4 2 2 ]   =   3 2 ' h d 6 f a 6 1 7 2 ;  
         r a m _ c e l l [           4 2 3 ]   =   3 2 ' h b 0 5 6 9 d 8 5 ;  
         r a m _ c e l l [           4 2 4 ]   =   3 2 ' h 7 6 d 2 e 2 3 3 ;  
         r a m _ c e l l [           4 2 5 ]   =   3 2 ' h 9 c 1 6 0 1 b a ;  
         r a m _ c e l l [           4 2 6 ]   =   3 2 ' h b 8 e 7 0 3 4 0 ;  
         r a m _ c e l l [           4 2 7 ]   =   3 2 ' h a d 5 4 a 4 d b ;  
         r a m _ c e l l [           4 2 8 ]   =   3 2 ' h c f f 8 f b 5 7 ;  
         r a m _ c e l l [           4 2 9 ]   =   3 2 ' h 1 0 3 c 2 6 6 6 ;  
         r a m _ c e l l [           4 3 0 ]   =   3 2 ' h 6 5 2 3 4 e 9 6 ;  
         r a m _ c e l l [           4 3 1 ]   =   3 2 ' h 1 9 9 f 2 9 8 e ;  
         r a m _ c e l l [           4 3 2 ]   =   3 2 ' h 3 b 8 d 7 e 1 2 ;  
         r a m _ c e l l [           4 3 3 ]   =   3 2 ' h 0 3 b 7 9 5 f f ;  
         r a m _ c e l l [           4 3 4 ]   =   3 2 ' h d 6 6 0 7 3 7 9 ;  
         r a m _ c e l l [           4 3 5 ]   =   3 2 ' h 9 e a d 4 3 c 6 ;  
         r a m _ c e l l [           4 3 6 ]   =   3 2 ' h 2 a 3 7 f 1 9 5 ;  
         r a m _ c e l l [           4 3 7 ]   =   3 2 ' h 5 6 0 9 b 8 9 3 ;  
         r a m _ c e l l [           4 3 8 ]   =   3 2 ' h b 0 8 a 7 2 4 5 ;  
         r a m _ c e l l [           4 3 9 ]   =   3 2 ' h c 1 7 8 b 9 9 3 ;  
         r a m _ c e l l [           4 4 0 ]   =   3 2 ' h d 7 d 2 7 2 1 2 ;  
         r a m _ c e l l [           4 4 1 ]   =   3 2 ' h b 5 4 5 a 5 e 4 ;  
         r a m _ c e l l [           4 4 2 ]   =   3 2 ' h 7 6 7 d c f 5 3 ;  
         r a m _ c e l l [           4 4 3 ]   =   3 2 ' h d f 1 6 d 2 d 8 ;  
         r a m _ c e l l [           4 4 4 ]   =   3 2 ' h 3 b 4 6 6 a 9 e ;  
         r a m _ c e l l [           4 4 5 ]   =   3 2 ' h 1 5 b e 1 4 2 7 ;  
         r a m _ c e l l [           4 4 6 ]   =   3 2 ' h b c 9 9 3 b f e ;  
         r a m _ c e l l [           4 4 7 ]   =   3 2 ' h 3 4 f 3 b 5 b e ;  
         r a m _ c e l l [           4 4 8 ]   =   3 2 ' h 1 3 1 4 b a 8 b ;  
         r a m _ c e l l [           4 4 9 ]   =   3 2 ' h 4 a 8 0 4 7 e f ;  
         r a m _ c e l l [           4 5 0 ]   =   3 2 ' h d 8 a 8 4 b f f ;  
         r a m _ c e l l [           4 5 1 ]   =   3 2 ' h 4 5 7 b c c e 1 ;  
         r a m _ c e l l [           4 5 2 ]   =   3 2 ' h c 2 c 6 f 3 8 3 ;  
         r a m _ c e l l [           4 5 3 ]   =   3 2 ' h 8 d 8 1 3 d b 0 ;  
         r a m _ c e l l [           4 5 4 ]   =   3 2 ' h 5 1 1 3 e 0 d 5 ;  
         r a m _ c e l l [           4 5 5 ]   =   3 2 ' h 9 8 f 2 f 4 2 b ;  
         r a m _ c e l l [           4 5 6 ]   =   3 2 ' h f 3 1 a 5 a 3 0 ;  
         r a m _ c e l l [           4 5 7 ]   =   3 2 ' h 7 f b 0 2 d 8 4 ;  
         r a m _ c e l l [           4 5 8 ]   =   3 2 ' h 5 d 6 d 8 d b 2 ;  
         r a m _ c e l l [           4 5 9 ]   =   3 2 ' h e 7 5 8 1 d e 7 ;  
         r a m _ c e l l [           4 6 0 ]   =   3 2 ' h 9 7 d 0 3 b f 3 ;  
         r a m _ c e l l [           4 6 1 ]   =   3 2 ' h b d f d d a c 7 ;  
         r a m _ c e l l [           4 6 2 ]   =   3 2 ' h 2 8 7 3 3 2 2 f ;  
         r a m _ c e l l [           4 6 3 ]   =   3 2 ' h 2 2 3 a 2 f 1 8 ;  
         r a m _ c e l l [           4 6 4 ]   =   3 2 ' h a f d b 1 5 d d ;  
         r a m _ c e l l [           4 6 5 ]   =   3 2 ' h 0 d b 8 3 9 5 d ;  
         r a m _ c e l l [           4 6 6 ]   =   3 2 ' h 3 9 2 4 f 2 7 6 ;  
         r a m _ c e l l [           4 6 7 ]   =   3 2 ' h 8 3 a e 6 c e 5 ;  
         r a m _ c e l l [           4 6 8 ]   =   3 2 ' h 3 5 1 0 a 6 2 9 ;  
         r a m _ c e l l [           4 6 9 ]   =   3 2 ' h a f c 7 f 6 4 d ;  
         r a m _ c e l l [           4 7 0 ]   =   3 2 ' h 2 3 b 3 0 9 5 4 ;  
         r a m _ c e l l [           4 7 1 ]   =   3 2 ' h 1 1 9 b e 1 c 0 ;  
         r a m _ c e l l [           4 7 2 ]   =   3 2 ' h e 8 7 9 9 1 c a ;  
         r a m _ c e l l [           4 7 3 ]   =   3 2 ' h d 9 1 2 0 8 3 a ;  
         r a m _ c e l l [           4 7 4 ]   =   3 2 ' h 1 4 8 1 4 c d b ;  
         r a m _ c e l l [           4 7 5 ]   =   3 2 ' h 5 d 8 6 5 a 9 8 ;  
         r a m _ c e l l [           4 7 6 ]   =   3 2 ' h d 2 5 3 f 9 7 5 ;  
         r a m _ c e l l [           4 7 7 ]   =   3 2 ' h 0 a f 0 4 2 f 4 ;  
         r a m _ c e l l [           4 7 8 ]   =   3 2 ' h 7 d 2 6 8 1 8 f ;  
         r a m _ c e l l [           4 7 9 ]   =   3 2 ' h c b e b 9 b c 6 ;  
         r a m _ c e l l [           4 8 0 ]   =   3 2 ' h 2 c 1 b 4 e c c ;  
         r a m _ c e l l [           4 8 1 ]   =   3 2 ' h 6 a 5 a 0 2 9 e ;  
         r a m _ c e l l [           4 8 2 ]   =   3 2 ' h 5 6 4 c 4 a c 4 ;  
         r a m _ c e l l [           4 8 3 ]   =   3 2 ' h 2 9 c 5 6 3 9 a ;  
         r a m _ c e l l [           4 8 4 ]   =   3 2 ' h 1 f f 8 3 3 6 6 ;  
         r a m _ c e l l [           4 8 5 ]   =   3 2 ' h 1 4 6 8 3 f 2 8 ;  
         r a m _ c e l l [           4 8 6 ]   =   3 2 ' h f 8 a d f 5 6 d ;  
         r a m _ c e l l [           4 8 7 ]   =   3 2 ' h 1 4 9 5 6 8 8 a ;  
         r a m _ c e l l [           4 8 8 ]   =   3 2 ' h 3 f 0 1 8 e 1 0 ;  
         r a m _ c e l l [           4 8 9 ]   =   3 2 ' h 3 4 f e c f 4 2 ;  
         r a m _ c e l l [           4 9 0 ]   =   3 2 ' h 3 2 2 d c 7 c 7 ;  
         r a m _ c e l l [           4 9 1 ]   =   3 2 ' h 4 6 f 7 1 8 2 d ;  
         r a m _ c e l l [           4 9 2 ]   =   3 2 ' h 0 f 7 d 5 b 9 f ;  
         r a m _ c e l l [           4 9 3 ]   =   3 2 ' h b 5 4 e b 1 4 2 ;  
         r a m _ c e l l [           4 9 4 ]   =   3 2 ' h d d f 6 6 4 0 b ;  
         r a m _ c e l l [           4 9 5 ]   =   3 2 ' h 8 3 a 7 8 0 6 9 ;  
         r a m _ c e l l [           4 9 6 ]   =   3 2 ' h c c 8 e b 4 4 8 ;  
         r a m _ c e l l [           4 9 7 ]   =   3 2 ' h c 3 4 a d a 7 7 ;  
         r a m _ c e l l [           4 9 8 ]   =   3 2 ' h 5 b f 9 b 3 a 2 ;  
         r a m _ c e l l [           4 9 9 ]   =   3 2 ' h a c 1 f 1 d 9 4 ;  
         r a m _ c e l l [           5 0 0 ]   =   3 2 ' h 2 3 f 3 5 c 6 e ;  
         r a m _ c e l l [           5 0 1 ]   =   3 2 ' h e 8 2 e 0 e c 1 ;  
         r a m _ c e l l [           5 0 2 ]   =   3 2 ' h 3 f c f 2 d e d ;  
         r a m _ c e l l [           5 0 3 ]   =   3 2 ' h 7 e a 3 2 5 b 0 ;  
         r a m _ c e l l [           5 0 4 ]   =   3 2 ' h c 1 f 5 9 c 7 3 ;  
         r a m _ c e l l [           5 0 5 ]   =   3 2 ' h 0 f 1 3 0 4 a 3 ;  
         r a m _ c e l l [           5 0 6 ]   =   3 2 ' h f 4 8 f 1 f c 6 ;  
         r a m _ c e l l [           5 0 7 ]   =   3 2 ' h e e 1 c a 8 a f ;  
         r a m _ c e l l [           5 0 8 ]   =   3 2 ' h 4 6 f 6 4 3 5 d ;  
         r a m _ c e l l [           5 0 9 ]   =   3 2 ' h 1 7 6 3 c 6 5 3 ;  
         r a m _ c e l l [           5 1 0 ]   =   3 2 ' h 3 4 e d c 0 6 7 ;  
         r a m _ c e l l [           5 1 1 ]   =   3 2 ' h 0 8 f f 1 1 b c ;  
         / /   s r c   m a t r i x   B  
         r a m _ c e l l [           5 1 2 ]   =   3 2 ' h b 6 2 a a d 3 c ;  
         r a m _ c e l l [           5 1 3 ]   =   3 2 ' h 5 1 d d 3 a a 1 ;  
         r a m _ c e l l [           5 1 4 ]   =   3 2 ' h 9 4 1 b 9 5 c 5 ;  
         r a m _ c e l l [           5 1 5 ]   =   3 2 ' h 1 7 e 3 e 9 b 1 ;  
         r a m _ c e l l [           5 1 6 ]   =   3 2 ' h 5 0 f 6 e 0 5 4 ;  
         r a m _ c e l l [           5 1 7 ]   =   3 2 ' h 9 d d 6 7 7 f 3 ;  
         r a m _ c e l l [           5 1 8 ]   =   3 2 ' h a d 4 6 9 9 5 4 ;  
         r a m _ c e l l [           5 1 9 ]   =   3 2 ' h 0 e 3 6 7 7 e 0 ;  
         r a m _ c e l l [           5 2 0 ]   =   3 2 ' h b 7 d 7 5 4 0 b ;  
         r a m _ c e l l [           5 2 1 ]   =   3 2 ' h 7 4 f d 8 1 7 9 ;  
         r a m _ c e l l [           5 2 2 ]   =   3 2 ' h a e 9 e c 2 d 8 ;  
         r a m _ c e l l [           5 2 3 ]   =   3 2 ' h f b f a 0 3 f 0 ;  
         r a m _ c e l l [           5 2 4 ]   =   3 2 ' h e 4 2 e 9 6 4 4 ;  
         r a m _ c e l l [           5 2 5 ]   =   3 2 ' h 7 9 1 c e 3 6 1 ;  
         r a m _ c e l l [           5 2 6 ]   =   3 2 ' h e 7 b 4 f 4 5 b ;  
         r a m _ c e l l [           5 2 7 ]   =   3 2 ' h 2 2 6 c 2 2 9 b ;  
         r a m _ c e l l [           5 2 8 ]   =   3 2 ' h e 3 7 b 4 a 2 0 ;  
         r a m _ c e l l [           5 2 9 ]   =   3 2 ' h 3 9 9 e 2 f 0 5 ;  
         r a m _ c e l l [           5 3 0 ]   =   3 2 ' h 3 f 8 9 6 0 f a ;  
         r a m _ c e l l [           5 3 1 ]   =   3 2 ' h f 1 4 0 f 7 3 8 ;  
         r a m _ c e l l [           5 3 2 ]   =   3 2 ' h 3 2 1 d a 7 5 e ;  
         r a m _ c e l l [           5 3 3 ]   =   3 2 ' h 6 0 2 f c e 7 f ;  
         r a m _ c e l l [           5 3 4 ]   =   3 2 ' h 0 1 4 d 3 5 1 9 ;  
         r a m _ c e l l [           5 3 5 ]   =   3 2 ' h 6 0 0 f 1 2 5 5 ;  
         r a m _ c e l l [           5 3 6 ]   =   3 2 ' h 4 5 0 c 0 b e a ;  
         r a m _ c e l l [           5 3 7 ]   =   3 2 ' h 8 e 1 0 b b c 0 ;  
         r a m _ c e l l [           5 3 8 ]   =   3 2 ' h 1 1 5 1 9 f d 6 ;  
         r a m _ c e l l [           5 3 9 ]   =   3 2 ' h b 2 2 6 e 9 8 5 ;  
         r a m _ c e l l [           5 4 0 ]   =   3 2 ' h 8 4 f 2 1 3 4 d ;  
         r a m _ c e l l [           5 4 1 ]   =   3 2 ' h 7 3 6 8 e 0 7 a ;  
         r a m _ c e l l [           5 4 2 ]   =   3 2 ' h 8 8 3 4 6 8 e e ;  
         r a m _ c e l l [           5 4 3 ]   =   3 2 ' h 4 c 8 4 8 a d d ;  
         r a m _ c e l l [           5 4 4 ]   =   3 2 ' h 7 5 3 5 0 3 4 a ;  
         r a m _ c e l l [           5 4 5 ]   =   3 2 ' h a b a b b 3 c f ;  
         r a m _ c e l l [           5 4 6 ]   =   3 2 ' h 2 f 4 d f a f 0 ;  
         r a m _ c e l l [           5 4 7 ]   =   3 2 ' h 2 3 c b f 2 f d ;  
         r a m _ c e l l [           5 4 8 ]   =   3 2 ' h 7 d f 8 b 1 0 9 ;  
         r a m _ c e l l [           5 4 9 ]   =   3 2 ' h 6 b 7 9 e f 6 a ;  
         r a m _ c e l l [           5 5 0 ]   =   3 2 ' h 6 a 5 b 1 8 4 c ;  
         r a m _ c e l l [           5 5 1 ]   =   3 2 ' h 1 c a e 2 9 4 5 ;  
         r a m _ c e l l [           5 5 2 ]   =   3 2 ' h c 0 8 8 f 4 7 a ;  
         r a m _ c e l l [           5 5 3 ]   =   3 2 ' h f 1 a 1 4 b 4 b ;  
         r a m _ c e l l [           5 5 4 ]   =   3 2 ' h a 4 b 0 6 6 9 7 ;  
         r a m _ c e l l [           5 5 5 ]   =   3 2 ' h 7 a c f d 8 f 9 ;  
         r a m _ c e l l [           5 5 6 ]   =   3 2 ' h b 2 a b b 4 0 2 ;  
         r a m _ c e l l [           5 5 7 ]   =   3 2 ' h e c c 6 0 c e 6 ;  
         r a m _ c e l l [           5 5 8 ]   =   3 2 ' h 5 e 7 5 e 5 c 9 ;  
         r a m _ c e l l [           5 5 9 ]   =   3 2 ' h 5 1 4 3 1 8 1 a ;  
         r a m _ c e l l [           5 6 0 ]   =   3 2 ' h 9 3 6 6 b f 7 e ;  
         r a m _ c e l l [           5 6 1 ]   =   3 2 ' h 5 e 9 2 9 f b 0 ;  
         r a m _ c e l l [           5 6 2 ]   =   3 2 ' h 0 2 0 0 1 5 c 9 ;  
         r a m _ c e l l [           5 6 3 ]   =   3 2 ' h d 7 5 f 4 6 b c ;  
         r a m _ c e l l [           5 6 4 ]   =   3 2 ' h b 7 d c 6 1 4 c ;  
         r a m _ c e l l [           5 6 5 ]   =   3 2 ' h 2 4 0 a 8 8 8 9 ;  
         r a m _ c e l l [           5 6 6 ]   =   3 2 ' h 9 7 b 0 8 8 0 3 ;  
         r a m _ c e l l [           5 6 7 ]   =   3 2 ' h 8 5 e c 3 8 9 9 ;  
         r a m _ c e l l [           5 6 8 ]   =   3 2 ' h e 5 d 7 4 b 8 b ;  
         r a m _ c e l l [           5 6 9 ]   =   3 2 ' h 5 4 5 5 1 3 d 3 ;  
         r a m _ c e l l [           5 7 0 ]   =   3 2 ' h 8 9 b a b 0 2 e ;  
         r a m _ c e l l [           5 7 1 ]   =   3 2 ' h 0 0 7 5 4 b b 8 ;  
         r a m _ c e l l [           5 7 2 ]   =   3 2 ' h 5 1 f 6 d 6 a 5 ;  
         r a m _ c e l l [           5 7 3 ]   =   3 2 ' h a 0 6 6 7 5 c 4 ;  
         r a m _ c e l l [           5 7 4 ]   =   3 2 ' h 9 3 e 0 7 c 3 9 ;  
         r a m _ c e l l [           5 7 5 ]   =   3 2 ' h d 0 d a f e 0 8 ;  
         r a m _ c e l l [           5 7 6 ]   =   3 2 ' h c b e e 5 4 9 d ;  
         r a m _ c e l l [           5 7 7 ]   =   3 2 ' h c a 4 1 a 5 9 8 ;  
         r a m _ c e l l [           5 7 8 ]   =   3 2 ' h f 2 e a c b 4 7 ;  
         r a m _ c e l l [           5 7 9 ]   =   3 2 ' h d 4 2 8 c 0 c 7 ;  
         r a m _ c e l l [           5 8 0 ]   =   3 2 ' h 9 a 9 0 d 2 3 4 ;  
         r a m _ c e l l [           5 8 1 ]   =   3 2 ' h e 4 1 7 5 d 7 3 ;  
         r a m _ c e l l [           5 8 2 ]   =   3 2 ' h 9 9 5 4 4 5 6 7 ;  
         r a m _ c e l l [           5 8 3 ]   =   3 2 ' h 6 2 0 8 b 4 d 9 ;  
         r a m _ c e l l [           5 8 4 ]   =   3 2 ' h 3 6 4 6 a d 2 d ;  
         r a m _ c e l l [           5 8 5 ]   =   3 2 ' h 3 2 4 b 2 d f e ;  
         r a m _ c e l l [           5 8 6 ]   =   3 2 ' h b 7 8 f d b 3 d ;  
         r a m _ c e l l [           5 8 7 ]   =   3 2 ' h d f 4 9 1 e e 3 ;  
         r a m _ c e l l [           5 8 8 ]   =   3 2 ' h 2 c 2 a 9 8 c 4 ;  
         r a m _ c e l l [           5 8 9 ]   =   3 2 ' h 2 9 d 1 d 7 8 9 ;  
         r a m _ c e l l [           5 9 0 ]   =   3 2 ' h b b c f 9 c a 3 ;  
         r a m _ c e l l [           5 9 1 ]   =   3 2 ' h 0 a b d 4 4 c e ;  
         r a m _ c e l l [           5 9 2 ]   =   3 2 ' h 9 6 a d a 6 7 1 ;  
         r a m _ c e l l [           5 9 3 ]   =   3 2 ' h 4 8 c f c 3 8 8 ;  
         r a m _ c e l l [           5 9 4 ]   =   3 2 ' h 3 2 0 b c 6 7 7 ;  
         r a m _ c e l l [           5 9 5 ]   =   3 2 ' h 3 c 3 a 5 c 4 8 ;  
         r a m _ c e l l [           5 9 6 ]   =   3 2 ' h d 1 a b f 4 d 5 ;  
         r a m _ c e l l [           5 9 7 ]   =   3 2 ' h 3 5 4 1 e 3 3 7 ;  
         r a m _ c e l l [           5 9 8 ]   =   3 2 ' h a 5 c 9 e c c d ;  
         r a m _ c e l l [           5 9 9 ]   =   3 2 ' h 7 a 5 e f 7 5 6 ;  
         r a m _ c e l l [           6 0 0 ]   =   3 2 ' h e 1 f f f a a 2 ;  
         r a m _ c e l l [           6 0 1 ]   =   3 2 ' h 3 d 8 4 e a 5 a ;  
         r a m _ c e l l [           6 0 2 ]   =   3 2 ' h 0 4 1 c 9 1 b 5 ;  
         r a m _ c e l l [           6 0 3 ]   =   3 2 ' h 3 8 d 9 7 b 2 9 ;  
         r a m _ c e l l [           6 0 4 ]   =   3 2 ' h 4 4 3 7 3 9 c 1 ;  
         r a m _ c e l l [           6 0 5 ]   =   3 2 ' h e 2 2 b 2 3 4 5 ;  
         r a m _ c e l l [           6 0 6 ]   =   3 2 ' h 8 e 6 5 9 a f 4 ;  
         r a m _ c e l l [           6 0 7 ]   =   3 2 ' h 7 c c 5 f 7 e b ;  
         r a m _ c e l l [           6 0 8 ]   =   3 2 ' h 2 c 5 f c 8 7 8 ;  
         r a m _ c e l l [           6 0 9 ]   =   3 2 ' h 2 0 e 9 3 5 3 0 ;  
         r a m _ c e l l [           6 1 0 ]   =   3 2 ' h e d 5 c 2 9 e d ;  
         r a m _ c e l l [           6 1 1 ]   =   3 2 ' h d a b 1 4 5 b 3 ;  
         r a m _ c e l l [           6 1 2 ]   =   3 2 ' h 3 7 7 a 3 2 a b ;  
         r a m _ c e l l [           6 1 3 ]   =   3 2 ' h f 6 5 8 d b b e ;  
         r a m _ c e l l [           6 1 4 ]   =   3 2 ' h d a 8 1 3 e f 1 ;  
         r a m _ c e l l [           6 1 5 ]   =   3 2 ' h 9 a 8 5 4 7 e 9 ;  
         r a m _ c e l l [           6 1 6 ]   =   3 2 ' h 2 c 7 9 9 2 5 3 ;  
         r a m _ c e l l [           6 1 7 ]   =   3 2 ' h 2 3 7 3 2 c 9 e ;  
         r a m _ c e l l [           6 1 8 ]   =   3 2 ' h 1 5 0 7 0 5 b 8 ;  
         r a m _ c e l l [           6 1 9 ]   =   3 2 ' h 0 3 0 d 3 a 9 b ;  
         r a m _ c e l l [           6 2 0 ]   =   3 2 ' h 9 0 0 1 e 9 7 a ;  
         r a m _ c e l l [           6 2 1 ]   =   3 2 ' h 6 5 f 0 4 c b 7 ;  
         r a m _ c e l l [           6 2 2 ]   =   3 2 ' h 0 8 a 6 b 4 c b ;  
         r a m _ c e l l [           6 2 3 ]   =   3 2 ' h 8 2 7 9 c b 7 f ;  
         r a m _ c e l l [           6 2 4 ]   =   3 2 ' h b a f 0 d 4 7 5 ;  
         r a m _ c e l l [           6 2 5 ]   =   3 2 ' h 7 5 5 d 3 4 0 f ;  
         r a m _ c e l l [           6 2 6 ]   =   3 2 ' h 5 f 2 4 6 7 8 c ;  
         r a m _ c e l l [           6 2 7 ]   =   3 2 ' h e a c 2 8 f 4 a ;  
         r a m _ c e l l [           6 2 8 ]   =   3 2 ' h 3 b 5 6 6 1 0 b ;  
         r a m _ c e l l [           6 2 9 ]   =   3 2 ' h f 4 e 7 9 4 5 4 ;  
         r a m _ c e l l [           6 3 0 ]   =   3 2 ' h 6 d 8 1 d 1 7 f ;  
         r a m _ c e l l [           6 3 1 ]   =   3 2 ' h b 6 9 0 d 7 2 1 ;  
         r a m _ c e l l [           6 3 2 ]   =   3 2 ' h 1 b c 1 b b 8 3 ;  
         r a m _ c e l l [           6 3 3 ]   =   3 2 ' h 9 9 9 e 4 3 c 5 ;  
         r a m _ c e l l [           6 3 4 ]   =   3 2 ' h 6 5 b f 4 b 5 2 ;  
         r a m _ c e l l [           6 3 5 ]   =   3 2 ' h 0 e 2 c 2 d e a ;  
         r a m _ c e l l [           6 3 6 ]   =   3 2 ' h b 9 6 5 0 8 3 1 ;  
         r a m _ c e l l [           6 3 7 ]   =   3 2 ' h 5 3 6 7 e d b 9 ;  
         r a m _ c e l l [           6 3 8 ]   =   3 2 ' h a c 0 1 b 7 f b ;  
         r a m _ c e l l [           6 3 9 ]   =   3 2 ' h 4 d b d 9 b b e ;  
         r a m _ c e l l [           6 4 0 ]   =   3 2 ' h 7 3 e a a 3 a 8 ;  
         r a m _ c e l l [           6 4 1 ]   =   3 2 ' h c a f a 5 6 a 7 ;  
         r a m _ c e l l [           6 4 2 ]   =   3 2 ' h 0 c 9 4 a 1 2 c ;  
         r a m _ c e l l [           6 4 3 ]   =   3 2 ' h 5 9 8 c c 3 f 9 ;  
         r a m _ c e l l [           6 4 4 ]   =   3 2 ' h f 1 2 5 2 1 6 8 ;  
         r a m _ c e l l [           6 4 5 ]   =   3 2 ' h 8 1 e 8 4 2 5 0 ;  
         r a m _ c e l l [           6 4 6 ]   =   3 2 ' h a b c f d b b 6 ;  
         r a m _ c e l l [           6 4 7 ]   =   3 2 ' h e 2 d 7 5 0 d 3 ;  
         r a m _ c e l l [           6 4 8 ]   =   3 2 ' h f 9 2 0 1 b e 2 ;  
         r a m _ c e l l [           6 4 9 ]   =   3 2 ' h 6 d 2 7 8 8 1 5 ;  
         r a m _ c e l l [           6 5 0 ]   =   3 2 ' h e c 6 5 0 4 b e ;  
         r a m _ c e l l [           6 5 1 ]   =   3 2 ' h d d 3 1 5 e e 1 ;  
         r a m _ c e l l [           6 5 2 ]   =   3 2 ' h 0 4 7 a a 2 6 5 ;  
         r a m _ c e l l [           6 5 3 ]   =   3 2 ' h 8 4 0 e 4 f 5 6 ;  
         r a m _ c e l l [           6 5 4 ]   =   3 2 ' h 2 c c 2 a d 4 9 ;  
         r a m _ c e l l [           6 5 5 ]   =   3 2 ' h 2 f 9 3 6 f 2 7 ;  
         r a m _ c e l l [           6 5 6 ]   =   3 2 ' h 3 3 e 8 4 6 7 2 ;  
         r a m _ c e l l [           6 5 7 ]   =   3 2 ' h 3 7 c 6 9 7 a 7 ;  
         r a m _ c e l l [           6 5 8 ]   =   3 2 ' h 1 6 a 8 2 8 0 5 ;  
         r a m _ c e l l [           6 5 9 ]   =   3 2 ' h d 5 0 5 c 0 4 e ;  
         r a m _ c e l l [           6 6 0 ]   =   3 2 ' h f f 1 d 4 c e b ;  
         r a m _ c e l l [           6 6 1 ]   =   3 2 ' h 8 f e 3 9 e e a ;  
         r a m _ c e l l [           6 6 2 ]   =   3 2 ' h 9 9 e 9 0 9 9 7 ;  
         r a m _ c e l l [           6 6 3 ]   =   3 2 ' h e 6 2 e a b 1 1 ;  
         r a m _ c e l l [           6 6 4 ]   =   3 2 ' h 0 3 4 9 6 3 7 c ;  
         r a m _ c e l l [           6 6 5 ]   =   3 2 ' h 9 1 b c 7 d f a ;  
         r a m _ c e l l [           6 6 6 ]   =   3 2 ' h b d 4 b 0 7 5 e ;  
         r a m _ c e l l [           6 6 7 ]   =   3 2 ' h 8 d 3 c f 7 1 5 ;  
         r a m _ c e l l [           6 6 8 ]   =   3 2 ' h 2 4 6 9 3 2 1 b ;  
         r a m _ c e l l [           6 6 9 ]   =   3 2 ' h f 8 d 9 9 4 a 0 ;  
         r a m _ c e l l [           6 7 0 ]   =   3 2 ' h 9 5 c f 9 c 6 5 ;  
         r a m _ c e l l [           6 7 1 ]   =   3 2 ' h 1 7 c 9 f a e 1 ;  
         r a m _ c e l l [           6 7 2 ]   =   3 2 ' h f 6 6 8 5 1 5 6 ;  
         r a m _ c e l l [           6 7 3 ]   =   3 2 ' h 8 c d 8 0 9 1 e ;  
         r a m _ c e l l [           6 7 4 ]   =   3 2 ' h 3 c c d b 6 7 a ;  
         r a m _ c e l l [           6 7 5 ]   =   3 2 ' h e 8 a e b 8 2 c ;  
         r a m _ c e l l [           6 7 6 ]   =   3 2 ' h 4 4 f 2 f f a 3 ;  
         r a m _ c e l l [           6 7 7 ]   =   3 2 ' h 1 3 3 b 3 a 3 5 ;  
         r a m _ c e l l [           6 7 8 ]   =   3 2 ' h 4 b 8 1 c 9 a 8 ;  
         r a m _ c e l l [           6 7 9 ]   =   3 2 ' h 9 f f 9 6 b e c ;  
         r a m _ c e l l [           6 8 0 ]   =   3 2 ' h b 6 9 a 5 2 0 1 ;  
         r a m _ c e l l [           6 8 1 ]   =   3 2 ' h c f f d 4 a 8 a ;  
         r a m _ c e l l [           6 8 2 ]   =   3 2 ' h e 4 2 1 0 e 8 c ;  
         r a m _ c e l l [           6 8 3 ]   =   3 2 ' h 5 a e 4 4 5 6 d ;  
         r a m _ c e l l [           6 8 4 ]   =   3 2 ' h 4 b a 9 3 9 9 8 ;  
         r a m _ c e l l [           6 8 5 ]   =   3 2 ' h 9 f 5 4 5 8 0 f ;  
         r a m _ c e l l [           6 8 6 ]   =   3 2 ' h b 6 9 5 0 d d 7 ;  
         r a m _ c e l l [           6 8 7 ]   =   3 2 ' h 7 6 e 7 4 1 c a ;  
         r a m _ c e l l [           6 8 8 ]   =   3 2 ' h e c 0 7 9 6 8 6 ;  
         r a m _ c e l l [           6 8 9 ]   =   3 2 ' h 4 b 1 1 1 6 c 1 ;  
         r a m _ c e l l [           6 9 0 ]   =   3 2 ' h d f 6 e a e 1 1 ;  
         r a m _ c e l l [           6 9 1 ]   =   3 2 ' h 2 8 9 f 8 c 4 4 ;  
         r a m _ c e l l [           6 9 2 ]   =   3 2 ' h e b b d 3 d c 9 ;  
         r a m _ c e l l [           6 9 3 ]   =   3 2 ' h 5 d 4 2 2 4 c a ;  
         r a m _ c e l l [           6 9 4 ]   =   3 2 ' h d 8 7 b 7 8 e 3 ;  
         r a m _ c e l l [           6 9 5 ]   =   3 2 ' h c 6 9 9 a 1 1 4 ;  
         r a m _ c e l l [           6 9 6 ]   =   3 2 ' h f 3 8 c 5 c f 2 ;  
         r a m _ c e l l [           6 9 7 ]   =   3 2 ' h 0 8 a e a 4 6 9 ;  
         r a m _ c e l l [           6 9 8 ]   =   3 2 ' h e 4 2 8 0 4 3 d ;  
         r a m _ c e l l [           6 9 9 ]   =   3 2 ' h 2 7 d d 6 0 f 2 ;  
         r a m _ c e l l [           7 0 0 ]   =   3 2 ' h 9 c b a 1 1 0 7 ;  
         r a m _ c e l l [           7 0 1 ]   =   3 2 ' h 6 d 0 b 2 2 2 b ;  
         r a m _ c e l l [           7 0 2 ]   =   3 2 ' h 0 e 4 5 f 0 8 d ;  
         r a m _ c e l l [           7 0 3 ]   =   3 2 ' h 4 9 4 a 9 e 7 4 ;  
         r a m _ c e l l [           7 0 4 ]   =   3 2 ' h d 0 7 1 a 2 b 2 ;  
         r a m _ c e l l [           7 0 5 ]   =   3 2 ' h d 7 a 1 2 3 7 7 ;  
         r a m _ c e l l [           7 0 6 ]   =   3 2 ' h 3 c 6 e 9 e 2 9 ;  
         r a m _ c e l l [           7 0 7 ]   =   3 2 ' h 8 9 6 9 7 6 9 6 ;  
         r a m _ c e l l [           7 0 8 ]   =   3 2 ' h b e f 6 2 7 0 1 ;  
         r a m _ c e l l [           7 0 9 ]   =   3 2 ' h 9 a 6 2 3 f 3 5 ;  
         r a m _ c e l l [           7 1 0 ]   =   3 2 ' h 2 f 5 f 2 3 4 c ;  
         r a m _ c e l l [           7 1 1 ]   =   3 2 ' h e b 9 e f 5 7 5 ;  
         r a m _ c e l l [           7 1 2 ]   =   3 2 ' h 0 b 5 0 8 3 2 3 ;  
         r a m _ c e l l [           7 1 3 ]   =   3 2 ' h f b 7 d 8 c e 2 ;  
         r a m _ c e l l [           7 1 4 ]   =   3 2 ' h a 9 e 7 8 6 7 7 ;  
         r a m _ c e l l [           7 1 5 ]   =   3 2 ' h 4 6 0 1 a 4 d 6 ;  
         r a m _ c e l l [           7 1 6 ]   =   3 2 ' h 2 1 a 9 d f 5 8 ;  
         r a m _ c e l l [           7 1 7 ]   =   3 2 ' h b 9 e f b 8 4 9 ;  
         r a m _ c e l l [           7 1 8 ]   =   3 2 ' h 5 7 9 c 5 1 c 1 ;  
         r a m _ c e l l [           7 1 9 ]   =   3 2 ' h 9 2 2 5 a e c 9 ;  
         r a m _ c e l l [           7 2 0 ]   =   3 2 ' h a c 5 2 7 8 2 0 ;  
         r a m _ c e l l [           7 2 1 ]   =   3 2 ' h 3 6 f a 5 5 2 1 ;  
         r a m _ c e l l [           7 2 2 ]   =   3 2 ' h 2 6 b b 5 3 9 9 ;  
         r a m _ c e l l [           7 2 3 ]   =   3 2 ' h f 3 c 9 e a b b ;  
         r a m _ c e l l [           7 2 4 ]   =   3 2 ' h 1 3 2 d 5 c b c ;  
         r a m _ c e l l [           7 2 5 ]   =   3 2 ' h 2 f c 7 f 2 7 0 ;  
         r a m _ c e l l [           7 2 6 ]   =   3 2 ' h b 8 8 1 d 5 c 7 ;  
         r a m _ c e l l [           7 2 7 ]   =   3 2 ' h 3 a 7 d 0 d c d ;  
         r a m _ c e l l [           7 2 8 ]   =   3 2 ' h a 9 f 3 6 2 d e ;  
         r a m _ c e l l [           7 2 9 ]   =   3 2 ' h 1 9 a 8 3 3 0 5 ;  
         r a m _ c e l l [           7 3 0 ]   =   3 2 ' h b f b b 0 3 c 5 ;  
         r a m _ c e l l [           7 3 1 ]   =   3 2 ' h 2 4 9 3 c d c f ;  
         r a m _ c e l l [           7 3 2 ]   =   3 2 ' h 9 3 3 7 9 1 1 9 ;  
         r a m _ c e l l [           7 3 3 ]   =   3 2 ' h 6 c 6 c 6 6 e 7 ;  
         r a m _ c e l l [           7 3 4 ]   =   3 2 ' h 7 a b 5 c 9 7 7 ;  
         r a m _ c e l l [           7 3 5 ]   =   3 2 ' h 3 1 d a 0 7 f 0 ;  
         r a m _ c e l l [           7 3 6 ]   =   3 2 ' h 3 2 4 f 5 1 b e ;  
         r a m _ c e l l [           7 3 7 ]   =   3 2 ' h e 7 f 8 d a d 7 ;  
         r a m _ c e l l [           7 3 8 ]   =   3 2 ' h 6 b 8 7 d 1 7 b ;  
         r a m _ c e l l [           7 3 9 ]   =   3 2 ' h 9 3 a 7 1 c e b ;  
         r a m _ c e l l [           7 4 0 ]   =   3 2 ' h 8 f 5 b 7 c b 6 ;  
         r a m _ c e l l [           7 4 1 ]   =   3 2 ' h c 7 8 6 1 7 1 a ;  
         r a m _ c e l l [           7 4 2 ]   =   3 2 ' h 7 3 d 3 b 9 0 9 ;  
         r a m _ c e l l [           7 4 3 ]   =   3 2 ' h 9 9 6 0 4 6 0 e ;  
         r a m _ c e l l [           7 4 4 ]   =   3 2 ' h 5 5 c 0 3 7 e b ;  
         r a m _ c e l l [           7 4 5 ]   =   3 2 ' h 1 0 6 b 6 f d 5 ;  
         r a m _ c e l l [           7 4 6 ]   =   3 2 ' h f 0 5 b 2 e 1 0 ;  
         r a m _ c e l l [           7 4 7 ]   =   3 2 ' h 4 9 2 8 f 8 7 2 ;  
         r a m _ c e l l [           7 4 8 ]   =   3 2 ' h 6 9 6 4 d 4 f e ;  
         r a m _ c e l l [           7 4 9 ]   =   3 2 ' h f e 5 d 4 0 3 0 ;  
         r a m _ c e l l [           7 5 0 ]   =   3 2 ' h c 0 7 7 1 f 9 3 ;  
         r a m _ c e l l [           7 5 1 ]   =   3 2 ' h 8 f e 0 7 0 5 c ;  
         r a m _ c e l l [           7 5 2 ]   =   3 2 ' h 8 2 c d 6 8 d a ;  
         r a m _ c e l l [           7 5 3 ]   =   3 2 ' h e 6 6 b d 1 5 e ;  
         r a m _ c e l l [           7 5 4 ]   =   3 2 ' h 3 4 5 1 3 d 7 a ;  
         r a m _ c e l l [           7 5 5 ]   =   3 2 ' h 2 2 e 4 5 2 6 d ;  
         r a m _ c e l l [           7 5 6 ]   =   3 2 ' h a 0 0 a 9 0 4 9 ;  
         r a m _ c e l l [           7 5 7 ]   =   3 2 ' h 1 1 d d 2 b 1 6 ;  
         r a m _ c e l l [           7 5 8 ]   =   3 2 ' h e 5 a b e 1 d 8 ;  
         r a m _ c e l l [           7 5 9 ]   =   3 2 ' h e 7 0 0 6 b e 6 ;  
         r a m _ c e l l [           7 6 0 ]   =   3 2 ' h 6 9 f f 1 2 2 c ;  
         r a m _ c e l l [           7 6 1 ]   =   3 2 ' h 7 5 4 e 9 9 f c ;  
         r a m _ c e l l [           7 6 2 ]   =   3 2 ' h 4 4 0 7 1 8 4 7 ;  
         r a m _ c e l l [           7 6 3 ]   =   3 2 ' h 2 d f f 6 b b b ;  
         r a m _ c e l l [           7 6 4 ]   =   3 2 ' h a 2 a e 9 7 9 e ;  
         r a m _ c e l l [           7 6 5 ]   =   3 2 ' h 1 0 5 8 0 e 1 e ;  
         r a m _ c e l l [           7 6 6 ]   =   3 2 ' h 2 8 d e 3 a f b ;  
         r a m _ c e l l [           7 6 7 ]   =   3 2 ' h 6 a 4 2 d 0 6 9 ;  
 e n d  
  
 e n d m o d u l e  
  
 