
module mem #(                   //
    parameter  ADDR_LEN  = 11   //
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req)
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h3b934201;
    ram_cell[       1] = 32'h0;  // 32'he662a3da;
    ram_cell[       2] = 32'h0;  // 32'h12a6fe40;
    ram_cell[       3] = 32'h0;  // 32'h35677fb2;
    ram_cell[       4] = 32'h0;  // 32'hd6e04585;
    ram_cell[       5] = 32'h0;  // 32'ha9a2f2b8;
    ram_cell[       6] = 32'h0;  // 32'h3782e34f;
    ram_cell[       7] = 32'h0;  // 32'h52808fc8;
    ram_cell[       8] = 32'h0;  // 32'h34f378da;
    ram_cell[       9] = 32'h0;  // 32'h45f62974;
    ram_cell[      10] = 32'h0;  // 32'h8eb22e52;
    ram_cell[      11] = 32'h0;  // 32'he8ed91d9;
    ram_cell[      12] = 32'h0;  // 32'hc5741862;
    ram_cell[      13] = 32'h0;  // 32'h621860e1;
    ram_cell[      14] = 32'h0;  // 32'h411d441c;
    ram_cell[      15] = 32'h0;  // 32'h8ca04603;
    ram_cell[      16] = 32'h0;  // 32'hd3cbac09;
    ram_cell[      17] = 32'h0;  // 32'h2e44694b;
    ram_cell[      18] = 32'h0;  // 32'hf995d5d9;
    ram_cell[      19] = 32'h0;  // 32'h852ec40b;
    ram_cell[      20] = 32'h0;  // 32'ha2e00095;
    ram_cell[      21] = 32'h0;  // 32'haf24c390;
    ram_cell[      22] = 32'h0;  // 32'h9e271bb0;
    ram_cell[      23] = 32'h0;  // 32'h29245d02;
    ram_cell[      24] = 32'h0;  // 32'hb4dcd47e;
    ram_cell[      25] = 32'h0;  // 32'he631cd3f;
    ram_cell[      26] = 32'h0;  // 32'hee19ca59;
    ram_cell[      27] = 32'h0;  // 32'h6918d224;
    ram_cell[      28] = 32'h0;  // 32'h1e644a80;
    ram_cell[      29] = 32'h0;  // 32'h467836a6;
    ram_cell[      30] = 32'h0;  // 32'hc167a22d;
    ram_cell[      31] = 32'h0;  // 32'h9a6978fc;
    ram_cell[      32] = 32'h0;  // 32'hf86e872c;
    ram_cell[      33] = 32'h0;  // 32'h599ed24f;
    ram_cell[      34] = 32'h0;  // 32'h2a6013c9;
    ram_cell[      35] = 32'h0;  // 32'h869d2098;
    ram_cell[      36] = 32'h0;  // 32'h49489195;
    ram_cell[      37] = 32'h0;  // 32'h341ac39d;
    ram_cell[      38] = 32'h0;  // 32'h0482c51a;
    ram_cell[      39] = 32'h0;  // 32'h426da1cd;
    ram_cell[      40] = 32'h0;  // 32'h06c2dc11;
    ram_cell[      41] = 32'h0;  // 32'haa0c12fd;
    ram_cell[      42] = 32'h0;  // 32'hb5ae47e8;
    ram_cell[      43] = 32'h0;  // 32'h1df3493b;
    ram_cell[      44] = 32'h0;  // 32'hf6b077c2;
    ram_cell[      45] = 32'h0;  // 32'heb2b1e7a;
    ram_cell[      46] = 32'h0;  // 32'h8f4ec471;
    ram_cell[      47] = 32'h0;  // 32'h8ea240b0;
    ram_cell[      48] = 32'h0;  // 32'he0c6805d;
    ram_cell[      49] = 32'h0;  // 32'h046e58d5;
    ram_cell[      50] = 32'h0;  // 32'h9520f40b;
    ram_cell[      51] = 32'h0;  // 32'hff56b055;
    ram_cell[      52] = 32'h0;  // 32'h32fcafff;
    ram_cell[      53] = 32'h0;  // 32'hd78108ed;
    ram_cell[      54] = 32'h0;  // 32'h6a81dcb4;
    ram_cell[      55] = 32'h0;  // 32'h7c38cc63;
    ram_cell[      56] = 32'h0;  // 32'h4e2f900c;
    ram_cell[      57] = 32'h0;  // 32'h781b0583;
    ram_cell[      58] = 32'h0;  // 32'h1c5d2afb;
    ram_cell[      59] = 32'h0;  // 32'hb1b254ab;
    ram_cell[      60] = 32'h0;  // 32'h76bfff68;
    ram_cell[      61] = 32'h0;  // 32'hf1d97f42;
    ram_cell[      62] = 32'h0;  // 32'h2ef407d4;
    ram_cell[      63] = 32'h0;  // 32'h7109140a;
    ram_cell[      64] = 32'h0;  // 32'h4474f5c5;
    ram_cell[      65] = 32'h0;  // 32'he64930c1;
    ram_cell[      66] = 32'h0;  // 32'h6eb5a1a4;
    ram_cell[      67] = 32'h0;  // 32'h5fb12e4f;
    ram_cell[      68] = 32'h0;  // 32'h28d3ce04;
    ram_cell[      69] = 32'h0;  // 32'h212e3ce8;
    ram_cell[      70] = 32'h0;  // 32'h0a9e258f;
    ram_cell[      71] = 32'h0;  // 32'h94d49f10;
    ram_cell[      72] = 32'h0;  // 32'h7e6a0d91;
    ram_cell[      73] = 32'h0;  // 32'he9382812;
    ram_cell[      74] = 32'h0;  // 32'h02198571;
    ram_cell[      75] = 32'h0;  // 32'hd78fb480;
    ram_cell[      76] = 32'h0;  // 32'h2569cb01;
    ram_cell[      77] = 32'h0;  // 32'h964ac8dc;
    ram_cell[      78] = 32'h0;  // 32'h6559255b;
    ram_cell[      79] = 32'h0;  // 32'hc4522bcb;
    ram_cell[      80] = 32'h0;  // 32'h7f452086;
    ram_cell[      81] = 32'h0;  // 32'h8762f594;
    ram_cell[      82] = 32'h0;  // 32'h7b68c226;
    ram_cell[      83] = 32'h0;  // 32'h5f537fbe;
    ram_cell[      84] = 32'h0;  // 32'h41116a20;
    ram_cell[      85] = 32'h0;  // 32'hb9f390d7;
    ram_cell[      86] = 32'h0;  // 32'hdf6c62e3;
    ram_cell[      87] = 32'h0;  // 32'h38d96a09;
    ram_cell[      88] = 32'h0;  // 32'h97f594d6;
    ram_cell[      89] = 32'h0;  // 32'h9c14390a;
    ram_cell[      90] = 32'h0;  // 32'hb0cd0b04;
    ram_cell[      91] = 32'h0;  // 32'h7f388c9c;
    ram_cell[      92] = 32'h0;  // 32'he069f59c;
    ram_cell[      93] = 32'h0;  // 32'hba246aac;
    ram_cell[      94] = 32'h0;  // 32'hd20d1c46;
    ram_cell[      95] = 32'h0;  // 32'h028d4c20;
    ram_cell[      96] = 32'h0;  // 32'h37e4b0ed;
    ram_cell[      97] = 32'h0;  // 32'hacad08a4;
    ram_cell[      98] = 32'h0;  // 32'he8075b5c;
    ram_cell[      99] = 32'h0;  // 32'h76ffd4ac;
    ram_cell[     100] = 32'h0;  // 32'hc7e8b755;
    ram_cell[     101] = 32'h0;  // 32'h16621ac9;
    ram_cell[     102] = 32'h0;  // 32'h78a7dd69;
    ram_cell[     103] = 32'h0;  // 32'ha8f14266;
    ram_cell[     104] = 32'h0;  // 32'hf4a579fc;
    ram_cell[     105] = 32'h0;  // 32'hc22699a5;
    ram_cell[     106] = 32'h0;  // 32'h3d405843;
    ram_cell[     107] = 32'h0;  // 32'h52c0d595;
    ram_cell[     108] = 32'h0;  // 32'h8d691e70;
    ram_cell[     109] = 32'h0;  // 32'h5f2d7bfe;
    ram_cell[     110] = 32'h0;  // 32'hda79b7ed;
    ram_cell[     111] = 32'h0;  // 32'hca2750e7;
    ram_cell[     112] = 32'h0;  // 32'h7c201720;
    ram_cell[     113] = 32'h0;  // 32'he5bf7608;
    ram_cell[     114] = 32'h0;  // 32'h2dd74ba8;
    ram_cell[     115] = 32'h0;  // 32'h53f7e506;
    ram_cell[     116] = 32'h0;  // 32'h85032a6b;
    ram_cell[     117] = 32'h0;  // 32'h02c5a68b;
    ram_cell[     118] = 32'h0;  // 32'h2462c078;
    ram_cell[     119] = 32'h0;  // 32'h55183e59;
    ram_cell[     120] = 32'h0;  // 32'h190d5b9f;
    ram_cell[     121] = 32'h0;  // 32'hd54826af;
    ram_cell[     122] = 32'h0;  // 32'h0f747c9e;
    ram_cell[     123] = 32'h0;  // 32'h6e99347e;
    ram_cell[     124] = 32'h0;  // 32'h6c88e614;
    ram_cell[     125] = 32'h0;  // 32'h96eb1c34;
    ram_cell[     126] = 32'h0;  // 32'h73811db3;
    ram_cell[     127] = 32'h0;  // 32'h33b49008;
    ram_cell[     128] = 32'h0;  // 32'h0e2370db;
    ram_cell[     129] = 32'h0;  // 32'h9ca92543;
    ram_cell[     130] = 32'h0;  // 32'h4e7c3267;
    ram_cell[     131] = 32'h0;  // 32'h7fa5637f;
    ram_cell[     132] = 32'h0;  // 32'he3d323c9;
    ram_cell[     133] = 32'h0;  // 32'hc821e6a1;
    ram_cell[     134] = 32'h0;  // 32'h3d3e74f4;
    ram_cell[     135] = 32'h0;  // 32'hcde1ff3c;
    ram_cell[     136] = 32'h0;  // 32'h6115b1d9;
    ram_cell[     137] = 32'h0;  // 32'ha785fe6b;
    ram_cell[     138] = 32'h0;  // 32'h09292257;
    ram_cell[     139] = 32'h0;  // 32'hc725aea9;
    ram_cell[     140] = 32'h0;  // 32'hf7598990;
    ram_cell[     141] = 32'h0;  // 32'hd48bb687;
    ram_cell[     142] = 32'h0;  // 32'h1239252d;
    ram_cell[     143] = 32'h0;  // 32'h34cd881f;
    ram_cell[     144] = 32'h0;  // 32'h782f1934;
    ram_cell[     145] = 32'h0;  // 32'h7a8b00ff;
    ram_cell[     146] = 32'h0;  // 32'ha13f7633;
    ram_cell[     147] = 32'h0;  // 32'h6cd9fdc8;
    ram_cell[     148] = 32'h0;  // 32'hb014d63d;
    ram_cell[     149] = 32'h0;  // 32'he9c14a06;
    ram_cell[     150] = 32'h0;  // 32'h1de24532;
    ram_cell[     151] = 32'h0;  // 32'h71c583cd;
    ram_cell[     152] = 32'h0;  // 32'ha47a639c;
    ram_cell[     153] = 32'h0;  // 32'h00068243;
    ram_cell[     154] = 32'h0;  // 32'h1792e653;
    ram_cell[     155] = 32'h0;  // 32'h2cd35f8b;
    ram_cell[     156] = 32'h0;  // 32'hf9494b83;
    ram_cell[     157] = 32'h0;  // 32'h329140b8;
    ram_cell[     158] = 32'h0;  // 32'hc5900ed8;
    ram_cell[     159] = 32'h0;  // 32'h64724fd8;
    ram_cell[     160] = 32'h0;  // 32'h83af7941;
    ram_cell[     161] = 32'h0;  // 32'h90d780dc;
    ram_cell[     162] = 32'h0;  // 32'h35d43a5e;
    ram_cell[     163] = 32'h0;  // 32'h622c5412;
    ram_cell[     164] = 32'h0;  // 32'h5a02f3cb;
    ram_cell[     165] = 32'h0;  // 32'h3f4a063e;
    ram_cell[     166] = 32'h0;  // 32'h4e0715f8;
    ram_cell[     167] = 32'h0;  // 32'hcdb4f4c1;
    ram_cell[     168] = 32'h0;  // 32'he8e77d7c;
    ram_cell[     169] = 32'h0;  // 32'ha03b0615;
    ram_cell[     170] = 32'h0;  // 32'h5e81ab6a;
    ram_cell[     171] = 32'h0;  // 32'h764b5b14;
    ram_cell[     172] = 32'h0;  // 32'h9aa10817;
    ram_cell[     173] = 32'h0;  // 32'h45ff52d8;
    ram_cell[     174] = 32'h0;  // 32'hd413c18c;
    ram_cell[     175] = 32'h0;  // 32'hc26fecfe;
    ram_cell[     176] = 32'h0;  // 32'he8b752f1;
    ram_cell[     177] = 32'h0;  // 32'h97e3cd84;
    ram_cell[     178] = 32'h0;  // 32'hf6d5b52a;
    ram_cell[     179] = 32'h0;  // 32'h2cabaa30;
    ram_cell[     180] = 32'h0;  // 32'h16132ef1;
    ram_cell[     181] = 32'h0;  // 32'h2fec71de;
    ram_cell[     182] = 32'h0;  // 32'ha09a6856;
    ram_cell[     183] = 32'h0;  // 32'h6215202a;
    ram_cell[     184] = 32'h0;  // 32'h1a2b3b86;
    ram_cell[     185] = 32'h0;  // 32'ha3a28a57;
    ram_cell[     186] = 32'h0;  // 32'h446ef454;
    ram_cell[     187] = 32'h0;  // 32'h9169b771;
    ram_cell[     188] = 32'h0;  // 32'hc2ae26ec;
    ram_cell[     189] = 32'h0;  // 32'hee0240f0;
    ram_cell[     190] = 32'h0;  // 32'h60023060;
    ram_cell[     191] = 32'h0;  // 32'hcf6d8785;
    ram_cell[     192] = 32'h0;  // 32'hc3cd51a4;
    ram_cell[     193] = 32'h0;  // 32'h1966c51a;
    ram_cell[     194] = 32'h0;  // 32'hb9dfcf58;
    ram_cell[     195] = 32'h0;  // 32'ha152fe44;
    ram_cell[     196] = 32'h0;  // 32'h055ed369;
    ram_cell[     197] = 32'h0;  // 32'hea73b9b1;
    ram_cell[     198] = 32'h0;  // 32'h72d7d734;
    ram_cell[     199] = 32'h0;  // 32'h5cd82bf6;
    ram_cell[     200] = 32'h0;  // 32'hae557907;
    ram_cell[     201] = 32'h0;  // 32'h65fa0273;
    ram_cell[     202] = 32'h0;  // 32'hc122b759;
    ram_cell[     203] = 32'h0;  // 32'hf2d52ff5;
    ram_cell[     204] = 32'h0;  // 32'h4dc003af;
    ram_cell[     205] = 32'h0;  // 32'h4fa82945;
    ram_cell[     206] = 32'h0;  // 32'hbbfac540;
    ram_cell[     207] = 32'h0;  // 32'hb120ae2e;
    ram_cell[     208] = 32'h0;  // 32'h70956dc8;
    ram_cell[     209] = 32'h0;  // 32'h950e1e2c;
    ram_cell[     210] = 32'h0;  // 32'h468eecc8;
    ram_cell[     211] = 32'h0;  // 32'ha91f17c7;
    ram_cell[     212] = 32'h0;  // 32'hac246a51;
    ram_cell[     213] = 32'h0;  // 32'h8d491143;
    ram_cell[     214] = 32'h0;  // 32'hec0dac1d;
    ram_cell[     215] = 32'h0;  // 32'ha73b2b1e;
    ram_cell[     216] = 32'h0;  // 32'h2f2e104c;
    ram_cell[     217] = 32'h0;  // 32'h26f6c459;
    ram_cell[     218] = 32'h0;  // 32'h917499a7;
    ram_cell[     219] = 32'h0;  // 32'h21d0e824;
    ram_cell[     220] = 32'h0;  // 32'h1f075a2f;
    ram_cell[     221] = 32'h0;  // 32'h963c6945;
    ram_cell[     222] = 32'h0;  // 32'h8ae7d628;
    ram_cell[     223] = 32'h0;  // 32'h71bba9a6;
    ram_cell[     224] = 32'h0;  // 32'h45f0f662;
    ram_cell[     225] = 32'h0;  // 32'h765ffe75;
    ram_cell[     226] = 32'h0;  // 32'h64895ec0;
    ram_cell[     227] = 32'h0;  // 32'h0606fad3;
    ram_cell[     228] = 32'h0;  // 32'hd7f39cdb;
    ram_cell[     229] = 32'h0;  // 32'h3e41fb12;
    ram_cell[     230] = 32'h0;  // 32'h7bde53cd;
    ram_cell[     231] = 32'h0;  // 32'h3804c3f0;
    ram_cell[     232] = 32'h0;  // 32'hc709cd3c;
    ram_cell[     233] = 32'h0;  // 32'h43eb367c;
    ram_cell[     234] = 32'h0;  // 32'hbd6952f5;
    ram_cell[     235] = 32'h0;  // 32'h7f513221;
    ram_cell[     236] = 32'h0;  // 32'h75f5c32d;
    ram_cell[     237] = 32'h0;  // 32'hfe73d9de;
    ram_cell[     238] = 32'h0;  // 32'h2228ea06;
    ram_cell[     239] = 32'h0;  // 32'hd6428ef1;
    ram_cell[     240] = 32'h0;  // 32'h9e430dff;
    ram_cell[     241] = 32'h0;  // 32'h514b95c5;
    ram_cell[     242] = 32'h0;  // 32'h95438edf;
    ram_cell[     243] = 32'h0;  // 32'h6f54b5bc;
    ram_cell[     244] = 32'h0;  // 32'h91e94f75;
    ram_cell[     245] = 32'h0;  // 32'h23081c73;
    ram_cell[     246] = 32'h0;  // 32'h5f364b89;
    ram_cell[     247] = 32'h0;  // 32'h4aa7e912;
    ram_cell[     248] = 32'h0;  // 32'h6f91997f;
    ram_cell[     249] = 32'h0;  // 32'h1569ff74;
    ram_cell[     250] = 32'h0;  // 32'h919cd808;
    ram_cell[     251] = 32'h0;  // 32'h79eea3fa;
    ram_cell[     252] = 32'h0;  // 32'h0563e4fe;
    ram_cell[     253] = 32'h0;  // 32'hb006cf61;
    ram_cell[     254] = 32'h0;  // 32'h29ab7c9d;
    ram_cell[     255] = 32'h0;  // 32'hb0b11c3a;
    // src matrix A
    ram_cell[     256] = 32'h112dbf53;
    ram_cell[     257] = 32'hfca89b6b;
    ram_cell[     258] = 32'h87d1821e;
    ram_cell[     259] = 32'h19b96823;
    ram_cell[     260] = 32'h3bc14bfc;
    ram_cell[     261] = 32'hdf2ef4d7;
    ram_cell[     262] = 32'h3c0413f0;
    ram_cell[     263] = 32'h4cc56a10;
    ram_cell[     264] = 32'hcaae7e97;
    ram_cell[     265] = 32'h766ba961;
    ram_cell[     266] = 32'hcf5d8499;
    ram_cell[     267] = 32'h04b484dc;
    ram_cell[     268] = 32'he9a4e2bb;
    ram_cell[     269] = 32'h7db97027;
    ram_cell[     270] = 32'h7253666a;
    ram_cell[     271] = 32'h65ad52cd;
    ram_cell[     272] = 32'h61dc573a;
    ram_cell[     273] = 32'hf96da03e;
    ram_cell[     274] = 32'h3a907c9a;
    ram_cell[     275] = 32'h6818dd9a;
    ram_cell[     276] = 32'h2fb16a27;
    ram_cell[     277] = 32'hf589524a;
    ram_cell[     278] = 32'h305a0c80;
    ram_cell[     279] = 32'h84458ac0;
    ram_cell[     280] = 32'h71005547;
    ram_cell[     281] = 32'h5f110e7f;
    ram_cell[     282] = 32'h80bd0cf2;
    ram_cell[     283] = 32'hf91a368c;
    ram_cell[     284] = 32'h4346e53b;
    ram_cell[     285] = 32'h81391392;
    ram_cell[     286] = 32'hbf779804;
    ram_cell[     287] = 32'hcff6e28f;
    ram_cell[     288] = 32'h10a60924;
    ram_cell[     289] = 32'h303e00ff;
    ram_cell[     290] = 32'h891ddd49;
    ram_cell[     291] = 32'hcb24c10f;
    ram_cell[     292] = 32'h76c6ea14;
    ram_cell[     293] = 32'h8ed2aa87;
    ram_cell[     294] = 32'h7ebeec6a;
    ram_cell[     295] = 32'hd3cf07b3;
    ram_cell[     296] = 32'h70017157;
    ram_cell[     297] = 32'he2919d15;
    ram_cell[     298] = 32'h50aa268f;
    ram_cell[     299] = 32'h3b287480;
    ram_cell[     300] = 32'h2dfa4735;
    ram_cell[     301] = 32'hd1c56546;
    ram_cell[     302] = 32'hb42edb47;
    ram_cell[     303] = 32'h796c7119;
    ram_cell[     304] = 32'h3af97341;
    ram_cell[     305] = 32'h079746aa;
    ram_cell[     306] = 32'h2384d319;
    ram_cell[     307] = 32'h0043e0b7;
    ram_cell[     308] = 32'hbbf5ab88;
    ram_cell[     309] = 32'hdfcb73a6;
    ram_cell[     310] = 32'ha1f4055f;
    ram_cell[     311] = 32'hb6e23fe1;
    ram_cell[     312] = 32'hc48c3d86;
    ram_cell[     313] = 32'h209061be;
    ram_cell[     314] = 32'he8e02c48;
    ram_cell[     315] = 32'h605b0478;
    ram_cell[     316] = 32'hfa2c2a8b;
    ram_cell[     317] = 32'h22e638ee;
    ram_cell[     318] = 32'h010c6b31;
    ram_cell[     319] = 32'h17eb54fb;
    ram_cell[     320] = 32'h932c0288;
    ram_cell[     321] = 32'h42a29d45;
    ram_cell[     322] = 32'h9a655f79;
    ram_cell[     323] = 32'hbaa89be5;
    ram_cell[     324] = 32'h216cf918;
    ram_cell[     325] = 32'hf1ab6617;
    ram_cell[     326] = 32'h1e60f5a8;
    ram_cell[     327] = 32'hbeba2b00;
    ram_cell[     328] = 32'h37c6e8d7;
    ram_cell[     329] = 32'h7e1f60d1;
    ram_cell[     330] = 32'hf3dc621f;
    ram_cell[     331] = 32'h8bf3adcd;
    ram_cell[     332] = 32'h07c057c8;
    ram_cell[     333] = 32'h8740985f;
    ram_cell[     334] = 32'hd44710fd;
    ram_cell[     335] = 32'h3433de3f;
    ram_cell[     336] = 32'h87fbf9b6;
    ram_cell[     337] = 32'ha80a204e;
    ram_cell[     338] = 32'hb2669ef0;
    ram_cell[     339] = 32'h9c62779c;
    ram_cell[     340] = 32'hdb058c8a;
    ram_cell[     341] = 32'h3b525b8a;
    ram_cell[     342] = 32'hd84f4baa;
    ram_cell[     343] = 32'had5d64ce;
    ram_cell[     344] = 32'hc020a116;
    ram_cell[     345] = 32'h318cd44d;
    ram_cell[     346] = 32'h378361c2;
    ram_cell[     347] = 32'h4960ea6e;
    ram_cell[     348] = 32'h8abf5599;
    ram_cell[     349] = 32'h4bc1f6c9;
    ram_cell[     350] = 32'h1ac37deb;
    ram_cell[     351] = 32'hf9bac460;
    ram_cell[     352] = 32'hedfed999;
    ram_cell[     353] = 32'h47fa887a;
    ram_cell[     354] = 32'hd8ab19a4;
    ram_cell[     355] = 32'h7f74654b;
    ram_cell[     356] = 32'h36d1f288;
    ram_cell[     357] = 32'h324f07dd;
    ram_cell[     358] = 32'h5e29c401;
    ram_cell[     359] = 32'h003aa470;
    ram_cell[     360] = 32'h2b69b765;
    ram_cell[     361] = 32'h350feef0;
    ram_cell[     362] = 32'he197f6c2;
    ram_cell[     363] = 32'hec6e92b6;
    ram_cell[     364] = 32'ha0a948fc;
    ram_cell[     365] = 32'h9870a549;
    ram_cell[     366] = 32'h6c7194cb;
    ram_cell[     367] = 32'h9bb9e4b1;
    ram_cell[     368] = 32'hb16f6c30;
    ram_cell[     369] = 32'h7e593b84;
    ram_cell[     370] = 32'h71d92c93;
    ram_cell[     371] = 32'hb7270c45;
    ram_cell[     372] = 32'h557ab441;
    ram_cell[     373] = 32'h7adc9ff3;
    ram_cell[     374] = 32'hd2572c82;
    ram_cell[     375] = 32'hec533bfe;
    ram_cell[     376] = 32'h7aa4edc4;
    ram_cell[     377] = 32'hfb03e044;
    ram_cell[     378] = 32'h77c4069e;
    ram_cell[     379] = 32'h20d13612;
    ram_cell[     380] = 32'ha4cde87c;
    ram_cell[     381] = 32'haa5f3d20;
    ram_cell[     382] = 32'h079a3b9b;
    ram_cell[     383] = 32'h56485227;
    ram_cell[     384] = 32'h20976319;
    ram_cell[     385] = 32'h01856203;
    ram_cell[     386] = 32'hbb3e2f73;
    ram_cell[     387] = 32'ha27eae8d;
    ram_cell[     388] = 32'hc34a26c6;
    ram_cell[     389] = 32'h4a7e10ab;
    ram_cell[     390] = 32'h3e707cb6;
    ram_cell[     391] = 32'h16bb65fc;
    ram_cell[     392] = 32'hf4402f50;
    ram_cell[     393] = 32'h4f50e119;
    ram_cell[     394] = 32'h19185332;
    ram_cell[     395] = 32'haff1944b;
    ram_cell[     396] = 32'hcfbaab31;
    ram_cell[     397] = 32'ha7f0500b;
    ram_cell[     398] = 32'h20d272be;
    ram_cell[     399] = 32'hdcd1523e;
    ram_cell[     400] = 32'hef1cc211;
    ram_cell[     401] = 32'hb7a940cb;
    ram_cell[     402] = 32'h86c47964;
    ram_cell[     403] = 32'h9918308e;
    ram_cell[     404] = 32'hc3a8b662;
    ram_cell[     405] = 32'h417a3f84;
    ram_cell[     406] = 32'hc3bdea69;
    ram_cell[     407] = 32'h2111683c;
    ram_cell[     408] = 32'h8e516c5c;
    ram_cell[     409] = 32'hcef393be;
    ram_cell[     410] = 32'h600b9153;
    ram_cell[     411] = 32'hfd0fc7ae;
    ram_cell[     412] = 32'h72edcf27;
    ram_cell[     413] = 32'h139239e0;
    ram_cell[     414] = 32'h139b14e4;
    ram_cell[     415] = 32'h176ef566;
    ram_cell[     416] = 32'h3a567bcb;
    ram_cell[     417] = 32'h9e8b00ff;
    ram_cell[     418] = 32'h4498a378;
    ram_cell[     419] = 32'h48a58e6b;
    ram_cell[     420] = 32'ha087b81e;
    ram_cell[     421] = 32'hff168f72;
    ram_cell[     422] = 32'hd6fa6172;
    ram_cell[     423] = 32'hb0569d85;
    ram_cell[     424] = 32'h76d2e233;
    ram_cell[     425] = 32'h9c1601ba;
    ram_cell[     426] = 32'hb8e70340;
    ram_cell[     427] = 32'had54a4db;
    ram_cell[     428] = 32'hcff8fb57;
    ram_cell[     429] = 32'h103c2666;
    ram_cell[     430] = 32'h65234e96;
    ram_cell[     431] = 32'h199f298e;
    ram_cell[     432] = 32'h3b8d7e12;
    ram_cell[     433] = 32'h03b795ff;
    ram_cell[     434] = 32'hd6607379;
    ram_cell[     435] = 32'h9ead43c6;
    ram_cell[     436] = 32'h2a37f195;
    ram_cell[     437] = 32'h5609b893;
    ram_cell[     438] = 32'hb08a7245;
    ram_cell[     439] = 32'hc178b993;
    ram_cell[     440] = 32'hd7d27212;
    ram_cell[     441] = 32'hb545a5e4;
    ram_cell[     442] = 32'h767dcf53;
    ram_cell[     443] = 32'hdf16d2d8;
    ram_cell[     444] = 32'h3b466a9e;
    ram_cell[     445] = 32'h15be1427;
    ram_cell[     446] = 32'hbc993bfe;
    ram_cell[     447] = 32'h34f3b5be;
    ram_cell[     448] = 32'h1314ba8b;
    ram_cell[     449] = 32'h4a8047ef;
    ram_cell[     450] = 32'hd8a84bff;
    ram_cell[     451] = 32'h457bcce1;
    ram_cell[     452] = 32'hc2c6f383;
    ram_cell[     453] = 32'h8d813db0;
    ram_cell[     454] = 32'h5113e0d5;
    ram_cell[     455] = 32'h98f2f42b;
    ram_cell[     456] = 32'hf31a5a30;
    ram_cell[     457] = 32'h7fb02d84;
    ram_cell[     458] = 32'h5d6d8db2;
    ram_cell[     459] = 32'he7581de7;
    ram_cell[     460] = 32'h97d03bf3;
    ram_cell[     461] = 32'hbdfddac7;
    ram_cell[     462] = 32'h2873322f;
    ram_cell[     463] = 32'h223a2f18;
    ram_cell[     464] = 32'hafdb15dd;
    ram_cell[     465] = 32'h0db8395d;
    ram_cell[     466] = 32'h3924f276;
    ram_cell[     467] = 32'h83ae6ce5;
    ram_cell[     468] = 32'h3510a629;
    ram_cell[     469] = 32'hafc7f64d;
    ram_cell[     470] = 32'h23b30954;
    ram_cell[     471] = 32'h119be1c0;
    ram_cell[     472] = 32'he87991ca;
    ram_cell[     473] = 32'hd912083a;
    ram_cell[     474] = 32'h14814cdb;
    ram_cell[     475] = 32'h5d865a98;
    ram_cell[     476] = 32'hd253f975;
    ram_cell[     477] = 32'h0af042f4;
    ram_cell[     478] = 32'h7d26818f;
    ram_cell[     479] = 32'hcbeb9bc6;
    ram_cell[     480] = 32'h2c1b4ecc;
    ram_cell[     481] = 32'h6a5a029e;
    ram_cell[     482] = 32'h564c4ac4;
    ram_cell[     483] = 32'h29c5639a;
    ram_cell[     484] = 32'h1ff83366;
    ram_cell[     485] = 32'h14683f28;
    ram_cell[     486] = 32'hf8adf56d;
    ram_cell[     487] = 32'h1495688a;
    ram_cell[     488] = 32'h3f018e10;
    ram_cell[     489] = 32'h34fecf42;
    ram_cell[     490] = 32'h322dc7c7;
    ram_cell[     491] = 32'h46f7182d;
    ram_cell[     492] = 32'h0f7d5b9f;
    ram_cell[     493] = 32'hb54eb142;
    ram_cell[     494] = 32'hddf6640b;
    ram_cell[     495] = 32'h83a78069;
    ram_cell[     496] = 32'hcc8eb448;
    ram_cell[     497] = 32'hc34ada77;
    ram_cell[     498] = 32'h5bf9b3a2;
    ram_cell[     499] = 32'hac1f1d94;
    ram_cell[     500] = 32'h23f35c6e;
    ram_cell[     501] = 32'he82e0ec1;
    ram_cell[     502] = 32'h3fcf2ded;
    ram_cell[     503] = 32'h7ea325b0;
    ram_cell[     504] = 32'hc1f59c73;
    ram_cell[     505] = 32'h0f1304a3;
    ram_cell[     506] = 32'hf48f1fc6;
    ram_cell[     507] = 32'hee1ca8af;
    ram_cell[     508] = 32'h46f6435d;
    ram_cell[     509] = 32'h1763c653;
    ram_cell[     510] = 32'h34edc067;
    ram_cell[     511] = 32'h08ff11bc;
    // src matrix B
    ram_cell[     512] = 32'hb62aad3c;
    ram_cell[     513] = 32'h51dd3aa1;
    ram_cell[     514] = 32'h941b95c5;
    ram_cell[     515] = 32'h17e3e9b1;
    ram_cell[     516] = 32'h50f6e054;
    ram_cell[     517] = 32'h9dd677f3;
    ram_cell[     518] = 32'had469954;
    ram_cell[     519] = 32'h0e3677e0;
    ram_cell[     520] = 32'hb7d7540b;
    ram_cell[     521] = 32'h74fd8179;
    ram_cell[     522] = 32'hae9ec2d8;
    ram_cell[     523] = 32'hfbfa03f0;
    ram_cell[     524] = 32'he42e9644;
    ram_cell[     525] = 32'h791ce361;
    ram_cell[     526] = 32'he7b4f45b;
    ram_cell[     527] = 32'h226c229b;
    ram_cell[     528] = 32'he37b4a20;
    ram_cell[     529] = 32'h399e2f05;
    ram_cell[     530] = 32'h3f8960fa;
    ram_cell[     531] = 32'hf140f738;
    ram_cell[     532] = 32'h321da75e;
    ram_cell[     533] = 32'h602fce7f;
    ram_cell[     534] = 32'h014d3519;
    ram_cell[     535] = 32'h600f1255;
    ram_cell[     536] = 32'h450c0bea;
    ram_cell[     537] = 32'h8e10bbc0;
    ram_cell[     538] = 32'h11519fd6;
    ram_cell[     539] = 32'hb226e985;
    ram_cell[     540] = 32'h84f2134d;
    ram_cell[     541] = 32'h7368e07a;
    ram_cell[     542] = 32'h883468ee;
    ram_cell[     543] = 32'h4c848add;
    ram_cell[     544] = 32'h7535034a;
    ram_cell[     545] = 32'hababb3cf;
    ram_cell[     546] = 32'h2f4dfaf0;
    ram_cell[     547] = 32'h23cbf2fd;
    ram_cell[     548] = 32'h7df8b109;
    ram_cell[     549] = 32'h6b79ef6a;
    ram_cell[     550] = 32'h6a5b184c;
    ram_cell[     551] = 32'h1cae2945;
    ram_cell[     552] = 32'hc088f47a;
    ram_cell[     553] = 32'hf1a14b4b;
    ram_cell[     554] = 32'ha4b06697;
    ram_cell[     555] = 32'h7acfd8f9;
    ram_cell[     556] = 32'hb2abb402;
    ram_cell[     557] = 32'hecc60ce6;
    ram_cell[     558] = 32'h5e75e5c9;
    ram_cell[     559] = 32'h5143181a;
    ram_cell[     560] = 32'h9366bf7e;
    ram_cell[     561] = 32'h5e929fb0;
    ram_cell[     562] = 32'h020015c9;
    ram_cell[     563] = 32'hd75f46bc;
    ram_cell[     564] = 32'hb7dc614c;
    ram_cell[     565] = 32'h240a8889;
    ram_cell[     566] = 32'h97b08803;
    ram_cell[     567] = 32'h85ec3899;
    ram_cell[     568] = 32'he5d74b8b;
    ram_cell[     569] = 32'h545513d3;
    ram_cell[     570] = 32'h89bab02e;
    ram_cell[     571] = 32'h00754bb8;
    ram_cell[     572] = 32'h51f6d6a5;
    ram_cell[     573] = 32'ha06675c4;
    ram_cell[     574] = 32'h93e07c39;
    ram_cell[     575] = 32'hd0dafe08;
    ram_cell[     576] = 32'hcbee549d;
    ram_cell[     577] = 32'hca41a598;
    ram_cell[     578] = 32'hf2eacb47;
    ram_cell[     579] = 32'hd428c0c7;
    ram_cell[     580] = 32'h9a90d234;
    ram_cell[     581] = 32'he4175d73;
    ram_cell[     582] = 32'h99544567;
    ram_cell[     583] = 32'h6208b4d9;
    ram_cell[     584] = 32'h3646ad2d;
    ram_cell[     585] = 32'h324b2dfe;
    ram_cell[     586] = 32'hb78fdb3d;
    ram_cell[     587] = 32'hdf491ee3;
    ram_cell[     588] = 32'h2c2a98c4;
    ram_cell[     589] = 32'h29d1d789;
    ram_cell[     590] = 32'hbbcf9ca3;
    ram_cell[     591] = 32'h0abd44ce;
    ram_cell[     592] = 32'h96ada671;
    ram_cell[     593] = 32'h48cfc388;
    ram_cell[     594] = 32'h320bc677;
    ram_cell[     595] = 32'h3c3a5c48;
    ram_cell[     596] = 32'hd1abf4d5;
    ram_cell[     597] = 32'h3541e337;
    ram_cell[     598] = 32'ha5c9eccd;
    ram_cell[     599] = 32'h7a5ef756;
    ram_cell[     600] = 32'he1fffaa2;
    ram_cell[     601] = 32'h3d84ea5a;
    ram_cell[     602] = 32'h041c91b5;
    ram_cell[     603] = 32'h38d97b29;
    ram_cell[     604] = 32'h443739c1;
    ram_cell[     605] = 32'he22b2345;
    ram_cell[     606] = 32'h8e659af4;
    ram_cell[     607] = 32'h7cc5f7eb;
    ram_cell[     608] = 32'h2c5fc878;
    ram_cell[     609] = 32'h20e93530;
    ram_cell[     610] = 32'hed5c29ed;
    ram_cell[     611] = 32'hdab145b3;
    ram_cell[     612] = 32'h377a32ab;
    ram_cell[     613] = 32'hf658dbbe;
    ram_cell[     614] = 32'hda813ef1;
    ram_cell[     615] = 32'h9a8547e9;
    ram_cell[     616] = 32'h2c799253;
    ram_cell[     617] = 32'h23732c9e;
    ram_cell[     618] = 32'h150705b8;
    ram_cell[     619] = 32'h030d3a9b;
    ram_cell[     620] = 32'h9001e97a;
    ram_cell[     621] = 32'h65f04cb7;
    ram_cell[     622] = 32'h08a6b4cb;
    ram_cell[     623] = 32'h8279cb7f;
    ram_cell[     624] = 32'hbaf0d475;
    ram_cell[     625] = 32'h755d340f;
    ram_cell[     626] = 32'h5f24678c;
    ram_cell[     627] = 32'heac28f4a;
    ram_cell[     628] = 32'h3b56610b;
    ram_cell[     629] = 32'hf4e79454;
    ram_cell[     630] = 32'h6d81d17f;
    ram_cell[     631] = 32'hb690d721;
    ram_cell[     632] = 32'h1bc1bb83;
    ram_cell[     633] = 32'h999e43c5;
    ram_cell[     634] = 32'h65bf4b52;
    ram_cell[     635] = 32'h0e2c2dea;
    ram_cell[     636] = 32'hb9650831;
    ram_cell[     637] = 32'h5367edb9;
    ram_cell[     638] = 32'hac01b7fb;
    ram_cell[     639] = 32'h4dbd9bbe;
    ram_cell[     640] = 32'h73eaa3a8;
    ram_cell[     641] = 32'hcafa56a7;
    ram_cell[     642] = 32'h0c94a12c;
    ram_cell[     643] = 32'h598cc3f9;
    ram_cell[     644] = 32'hf1252168;
    ram_cell[     645] = 32'h81e84250;
    ram_cell[     646] = 32'habcfdbb6;
    ram_cell[     647] = 32'he2d750d3;
    ram_cell[     648] = 32'hf9201be2;
    ram_cell[     649] = 32'h6d278815;
    ram_cell[     650] = 32'hec6504be;
    ram_cell[     651] = 32'hdd315ee1;
    ram_cell[     652] = 32'h047aa265;
    ram_cell[     653] = 32'h840e4f56;
    ram_cell[     654] = 32'h2cc2ad49;
    ram_cell[     655] = 32'h2f936f27;
    ram_cell[     656] = 32'h33e84672;
    ram_cell[     657] = 32'h37c697a7;
    ram_cell[     658] = 32'h16a82805;
    ram_cell[     659] = 32'hd505c04e;
    ram_cell[     660] = 32'hff1d4ceb;
    ram_cell[     661] = 32'h8fe39eea;
    ram_cell[     662] = 32'h99e90997;
    ram_cell[     663] = 32'he62eab11;
    ram_cell[     664] = 32'h0349637c;
    ram_cell[     665] = 32'h91bc7dfa;
    ram_cell[     666] = 32'hbd4b075e;
    ram_cell[     667] = 32'h8d3cf715;
    ram_cell[     668] = 32'h2469321b;
    ram_cell[     669] = 32'hf8d994a0;
    ram_cell[     670] = 32'h95cf9c65;
    ram_cell[     671] = 32'h17c9fae1;
    ram_cell[     672] = 32'hf6685156;
    ram_cell[     673] = 32'h8cd8091e;
    ram_cell[     674] = 32'h3ccdb67a;
    ram_cell[     675] = 32'he8aeb82c;
    ram_cell[     676] = 32'h44f2ffa3;
    ram_cell[     677] = 32'h133b3a35;
    ram_cell[     678] = 32'h4b81c9a8;
    ram_cell[     679] = 32'h9ff96bec;
    ram_cell[     680] = 32'hb69a5201;
    ram_cell[     681] = 32'hcffd4a8a;
    ram_cell[     682] = 32'he4210e8c;
    ram_cell[     683] = 32'h5ae4456d;
    ram_cell[     684] = 32'h4ba93998;
    ram_cell[     685] = 32'h9f54580f;
    ram_cell[     686] = 32'hb6950dd7;
    ram_cell[     687] = 32'h76e741ca;
    ram_cell[     688] = 32'hec079686;
    ram_cell[     689] = 32'h4b1116c1;
    ram_cell[     690] = 32'hdf6eae11;
    ram_cell[     691] = 32'h289f8c44;
    ram_cell[     692] = 32'hebbd3dc9;
    ram_cell[     693] = 32'h5d4224ca;
    ram_cell[     694] = 32'hd87b78e3;
    ram_cell[     695] = 32'hc699a114;
    ram_cell[     696] = 32'hf38c5cf2;
    ram_cell[     697] = 32'h08aea469;
    ram_cell[     698] = 32'he428043d;
    ram_cell[     699] = 32'h27dd60f2;
    ram_cell[     700] = 32'h9cba1107;
    ram_cell[     701] = 32'h6d0b222b;
    ram_cell[     702] = 32'h0e45f08d;
    ram_cell[     703] = 32'h494a9e74;
    ram_cell[     704] = 32'hd071a2b2;
    ram_cell[     705] = 32'hd7a12377;
    ram_cell[     706] = 32'h3c6e9e29;
    ram_cell[     707] = 32'h89697696;
    ram_cell[     708] = 32'hbef62701;
    ram_cell[     709] = 32'h9a623f35;
    ram_cell[     710] = 32'h2f5f234c;
    ram_cell[     711] = 32'heb9ef575;
    ram_cell[     712] = 32'h0b508323;
    ram_cell[     713] = 32'hfb7d8ce2;
    ram_cell[     714] = 32'ha9e78677;
    ram_cell[     715] = 32'h4601a4d6;
    ram_cell[     716] = 32'h21a9df58;
    ram_cell[     717] = 32'hb9efb849;
    ram_cell[     718] = 32'h579c51c1;
    ram_cell[     719] = 32'h9225aec9;
    ram_cell[     720] = 32'hac527820;
    ram_cell[     721] = 32'h36fa5521;
    ram_cell[     722] = 32'h26bb5399;
    ram_cell[     723] = 32'hf3c9eabb;
    ram_cell[     724] = 32'h132d5cbc;
    ram_cell[     725] = 32'h2fc7f270;
    ram_cell[     726] = 32'hb881d5c7;
    ram_cell[     727] = 32'h3a7d0dcd;
    ram_cell[     728] = 32'ha9f362de;
    ram_cell[     729] = 32'h19a83305;
    ram_cell[     730] = 32'hbfbb03c5;
    ram_cell[     731] = 32'h2493cdcf;
    ram_cell[     732] = 32'h93379119;
    ram_cell[     733] = 32'h6c6c66e7;
    ram_cell[     734] = 32'h7ab5c977;
    ram_cell[     735] = 32'h31da07f0;
    ram_cell[     736] = 32'h324f51be;
    ram_cell[     737] = 32'he7f8dad7;
    ram_cell[     738] = 32'h6b87d17b;
    ram_cell[     739] = 32'h93a71ceb;
    ram_cell[     740] = 32'h8f5b7cb6;
    ram_cell[     741] = 32'hc786171a;
    ram_cell[     742] = 32'h73d3b909;
    ram_cell[     743] = 32'h9960460e;
    ram_cell[     744] = 32'h55c037eb;
    ram_cell[     745] = 32'h106b6fd5;
    ram_cell[     746] = 32'hf05b2e10;
    ram_cell[     747] = 32'h4928f872;
    ram_cell[     748] = 32'h6964d4fe;
    ram_cell[     749] = 32'hfe5d4030;
    ram_cell[     750] = 32'hc0771f93;
    ram_cell[     751] = 32'h8fe0705c;
    ram_cell[     752] = 32'h82cd68da;
    ram_cell[     753] = 32'he66bd15e;
    ram_cell[     754] = 32'h34513d7a;
    ram_cell[     755] = 32'h22e4526d;
    ram_cell[     756] = 32'ha00a9049;
    ram_cell[     757] = 32'h11dd2b16;
    ram_cell[     758] = 32'he5abe1d8;
    ram_cell[     759] = 32'he7006be6;
    ram_cell[     760] = 32'h69ff122c;
    ram_cell[     761] = 32'h754e99fc;
    ram_cell[     762] = 32'h44071847;
    ram_cell[     763] = 32'h2dff6bbb;
    ram_cell[     764] = 32'ha2ae979e;
    ram_cell[     765] = 32'h10580e1e;
    ram_cell[     766] = 32'h28de3afb;
    ram_cell[     767] = 32'h6a42d069;
end

endmodule

